library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.regionizer_data.all;

entity regionizer_nomerge is
    port(
            ap_clk : IN STD_LOGIC;
            ap_rst : IN STD_LOGIC;
            ap_start : IN STD_LOGIC;
            ap_done : OUT STD_LOGIC;
            ap_idle : OUT STD_LOGIC;
            ap_ready : OUT STD_LOGIC;
            newevent : IN STD_LOGIC;
            tracks_in_0_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_3_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_3_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_4_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_4_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_5_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_5_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_6_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_6_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_7_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_7_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_8_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_8_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_0_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_3_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_3_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_4_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_4_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_5_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_5_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_6_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_6_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_7_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_7_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_8_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_8_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_0_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_0_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_0_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_0_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_0_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_0_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_1_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_1_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_1_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_1_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_1_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_1_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_2_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_2_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_2_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_2_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_2_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_2_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_3_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_3_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_3_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_3_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_3_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_3_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_4_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_4_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_4_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_4_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_4_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_4_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_5_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_5_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_5_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_5_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_5_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_5_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_6_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_6_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_6_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_6_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_6_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_6_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_7_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_7_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_7_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_7_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_7_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_7_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_8_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_8_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_8_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_8_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_8_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_8_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_9_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_9_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_9_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_9_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_9_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_9_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_9_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_9_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_10_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_10_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_10_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_10_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_10_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_10_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_10_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_10_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_11_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_11_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_11_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_11_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_11_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_11_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_11_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_11_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_12_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_12_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_12_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_12_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_12_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_12_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_12_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_12_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_13_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_13_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_13_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_13_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_13_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_13_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_13_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_13_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_14_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_14_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_14_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_14_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_14_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_14_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_14_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_14_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_15_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_15_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_15_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_15_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_15_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_15_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_15_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_15_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_16_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_16_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_16_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_16_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_16_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_16_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_16_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_16_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_17_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_17_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_17_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_17_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_17_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_17_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_17_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_17_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_18_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_18_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_18_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_18_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_18_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_18_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_18_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_18_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_19_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_19_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_19_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_19_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_19_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_19_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_19_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_19_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_20_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_20_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_20_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_20_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_20_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_20_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_20_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_20_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_21_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_21_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_21_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_21_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_21_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_21_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_21_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_21_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_22_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_22_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_22_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_22_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_22_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_22_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_22_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_22_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_23_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_23_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_23_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_23_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_23_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_23_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_23_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_23_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_24_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_24_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_24_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_24_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_24_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_24_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_24_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_24_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_25_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_25_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_25_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_25_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_25_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_25_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_25_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_25_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_26_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_26_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_26_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_26_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_26_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_26_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_26_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_26_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_27_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_27_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_27_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_27_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_27_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_27_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_27_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_27_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_28_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_28_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_28_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_28_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_28_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_28_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_28_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_28_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_29_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_29_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_29_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_29_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_29_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_29_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_29_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_29_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_30_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_30_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_30_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_30_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_30_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_30_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_30_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_30_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_31_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_31_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_31_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_31_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_31_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_31_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_31_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_31_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_32_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_32_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_32_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_32_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_32_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_32_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_32_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_32_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_33_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_33_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_33_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_33_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_33_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_33_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_33_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_33_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_34_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_34_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_34_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_34_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_34_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_34_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_34_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_34_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_35_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_35_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_35_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_35_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_35_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_35_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_35_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_35_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_36_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_36_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_36_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_36_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_36_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_36_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_36_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_36_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_37_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_37_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_37_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_37_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_37_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_37_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_37_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_37_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_38_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_38_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_38_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_38_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_38_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_38_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_38_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_38_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_39_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_39_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_39_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_39_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_39_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_39_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_39_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_39_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_40_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_40_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_40_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_40_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_40_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_40_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_40_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_40_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_41_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_41_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_41_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_41_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_41_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_41_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_41_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_41_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_42_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_42_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_42_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_42_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_42_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_42_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_42_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_42_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_43_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_43_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_43_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_43_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_43_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_43_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_43_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_43_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_44_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_44_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_44_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_44_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_44_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_44_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_44_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_44_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_45_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_45_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_45_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_45_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_45_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_45_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_45_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_45_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_46_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_46_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_46_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_46_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_46_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_46_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_46_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_46_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_47_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_47_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_47_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_47_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_47_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_47_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_47_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_47_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_48_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_48_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_48_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_48_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_48_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_48_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_48_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_48_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_49_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_49_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_49_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_49_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_49_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_49_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_49_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_49_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_50_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_50_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_50_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_50_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_50_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_50_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_50_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_50_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_51_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_51_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_51_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_51_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_51_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_51_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_51_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_51_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_52_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_52_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_52_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_52_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_52_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_52_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_52_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_52_rest_V_ap_vld : OUT STD_LOGIC;
            tracks_out_53_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_53_pt_V_ap_vld : OUT STD_LOGIC;
            tracks_out_53_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_53_eta_V_ap_vld : OUT STD_LOGIC;
            tracks_out_53_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_53_phi_V_ap_vld : OUT STD_LOGIC;
            tracks_out_53_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_53_rest_V_ap_vld : OUT STD_LOGIC;
            newevent_out : OUT STD_LOGIC;
            newevent_out_ap_vld : OUT STD_LOGIC 
    );
end regionizer_nomerge;

architecture Behavioral of regionizer_nomerge is
    constant NREGIONS : natural := NSECTORS*NFIFOS;

    signal links_in :       particles(NSECTORS*NFIBERS-1 downto 0);
    signal fifo_in :        particles(NREGIONS-1 downto 0);
    signal fifo_in_write :  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal fifo_in_roll  :  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');

    signal fifo_out :        particles(NREGIONS-1 downto 0);
    signal fifo_out_valid :  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal fifo_out_roll:    std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal regions_out :      particles(NREGIONS-1 downto 0);
    signal regions_out_valid: std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal regions_out_roll:  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');

begin

    gen_fifos: for ireg in NREGIONS-1 downto 0 generate
        reg_buffer : entity work.rolling_fifo
                        --generic map(FIFO_INDEX => ireg+1)
                        port map(ap_clk => ap_clk, 
                                 d_in    => fifo_in(ireg),
                                 write_in  => fifo_in_write(ireg),
                                 roll   => fifo_in_roll(ireg),
                                 d_out    => fifo_out(ireg),
                                 valid_out  => fifo_out_valid(ireg),
                                 full  => '0',
                                 roll_out  => fifo_out_roll(ireg)
                             );
    end generate;
   
    links_in( 0).pt <= unsigned(tracks_in_0_0_pt_V);
    links_in( 1).pt <= unsigned(tracks_in_0_1_pt_V);
    links_in( 2).pt <= unsigned(tracks_in_1_0_pt_V);
    links_in( 3).pt <= unsigned(tracks_in_1_1_pt_V);
    links_in( 4).pt <= unsigned(tracks_in_2_0_pt_V);
    links_in( 5).pt <= unsigned(tracks_in_2_1_pt_V);
    links_in( 6).pt <= unsigned(tracks_in_3_0_pt_V);
    links_in( 7).pt <= unsigned(tracks_in_3_1_pt_V);
    links_in( 8).pt <= unsigned(tracks_in_4_0_pt_V);
    links_in( 9).pt <= unsigned(tracks_in_4_1_pt_V);
    links_in(10).pt <= unsigned(tracks_in_5_0_pt_V);
    links_in(11).pt <= unsigned(tracks_in_5_1_pt_V);
    links_in(12).pt <= unsigned(tracks_in_6_0_pt_V);
    links_in(13).pt <= unsigned(tracks_in_6_1_pt_V);
    links_in(14).pt <= unsigned(tracks_in_7_0_pt_V);
    links_in(15).pt <= unsigned(tracks_in_7_1_pt_V);
    links_in(16).pt <= unsigned(tracks_in_8_0_pt_V);
    links_in(17).pt <= unsigned(tracks_in_8_1_pt_V);
    links_in( 0).eta <= signed(tracks_in_0_0_eta_V);
    links_in( 1).eta <= signed(tracks_in_0_1_eta_V);
    links_in( 2).eta <= signed(tracks_in_1_0_eta_V);
    links_in( 3).eta <= signed(tracks_in_1_1_eta_V);
    links_in( 4).eta <= signed(tracks_in_2_0_eta_V);
    links_in( 5).eta <= signed(tracks_in_2_1_eta_V);
    links_in( 6).eta <= signed(tracks_in_3_0_eta_V);
    links_in( 7).eta <= signed(tracks_in_3_1_eta_V);
    links_in( 8).eta <= signed(tracks_in_4_0_eta_V);
    links_in( 9).eta <= signed(tracks_in_4_1_eta_V);
    links_in(10).eta <= signed(tracks_in_5_0_eta_V);
    links_in(11).eta <= signed(tracks_in_5_1_eta_V);
    links_in(12).eta <= signed(tracks_in_6_0_eta_V);
    links_in(13).eta <= signed(tracks_in_6_1_eta_V);
    links_in(14).eta <= signed(tracks_in_7_0_eta_V);
    links_in(15).eta <= signed(tracks_in_7_1_eta_V);
    links_in(16).eta <= signed(tracks_in_8_0_eta_V);
    links_in(17).eta <= signed(tracks_in_8_1_eta_V);
    links_in( 0).phi <= signed(tracks_in_0_0_phi_V);
    links_in( 1).phi <= signed(tracks_in_0_1_phi_V);
    links_in( 2).phi <= signed(tracks_in_1_0_phi_V);
    links_in( 3).phi <= signed(tracks_in_1_1_phi_V);
    links_in( 4).phi <= signed(tracks_in_2_0_phi_V);
    links_in( 5).phi <= signed(tracks_in_2_1_phi_V);
    links_in( 6).phi <= signed(tracks_in_3_0_phi_V);
    links_in( 7).phi <= signed(tracks_in_3_1_phi_V);
    links_in( 8).phi <= signed(tracks_in_4_0_phi_V);
    links_in( 9).phi <= signed(tracks_in_4_1_phi_V);
    links_in(10).phi <= signed(tracks_in_5_0_phi_V);
    links_in(11).phi <= signed(tracks_in_5_1_phi_V);
    links_in(12).phi <= signed(tracks_in_6_0_phi_V);
    links_in(13).phi <= signed(tracks_in_6_1_phi_V);
    links_in(14).phi <= signed(tracks_in_7_0_phi_V);
    links_in(15).phi <= signed(tracks_in_7_1_phi_V);
    links_in(16).phi <= signed(tracks_in_8_0_phi_V);
    links_in(17).phi <= signed(tracks_in_8_1_phi_V);
    links_in( 0).rest <= unsigned(tracks_in_0_0_rest_V);
    links_in( 1).rest <= unsigned(tracks_in_0_1_rest_V);
    links_in( 2).rest <= unsigned(tracks_in_1_0_rest_V);
    links_in( 3).rest <= unsigned(tracks_in_1_1_rest_V);
    links_in( 4).rest <= unsigned(tracks_in_2_0_rest_V);
    links_in( 5).rest <= unsigned(tracks_in_2_1_rest_V);
    links_in( 6).rest <= unsigned(tracks_in_3_0_rest_V);
    links_in( 7).rest <= unsigned(tracks_in_3_1_rest_V);
    links_in( 8).rest <= unsigned(tracks_in_4_0_rest_V);
    links_in( 9).rest <= unsigned(tracks_in_4_1_rest_V);
    links_in(10).rest <= unsigned(tracks_in_5_0_rest_V);
    links_in(11).rest <= unsigned(tracks_in_5_1_rest_V);
    links_in(12).rest <= unsigned(tracks_in_6_0_rest_V);
    links_in(13).rest <= unsigned(tracks_in_6_1_rest_V);
    links_in(14).rest <= unsigned(tracks_in_7_0_rest_V);
    links_in(15).rest <= unsigned(tracks_in_7_1_rest_V);
    links_in(16).rest <= unsigned(tracks_in_8_0_rest_V);
    links_in(17).rest <= unsigned(tracks_in_8_1_rest_V);


    link2fifo : process(ap_clk)
        variable isec_next, isec_prev : integer range 0 to NSECTORS-1;
        variable link_this, link_next, link_prev : std_logic;
    begin
        if rising_edge(ap_clk) then
            for isec in 0 to NSECTORS-1 loop
                if isec = 0 then
                    isec_next := isec + 1;
                    isec_prev := NSECTORS-1;
                elsif isec = NSECTORS-1 then
                    isec_next := 0;
                    isec_prev := isec - 1;
                else
                    isec_next := isec + 1;
                    isec_prev := isec - 1;
                end if;
                for ifib in 0 to NFIBERS-1 loop
                    if ap_start = '0' or links_in(isec*NFIBERS+ifib).pt = 0 then
                        link_this := '0';
                        link_prev := '0';
                        link_next := '0';
                    else
                        link_this := '1';
                        if links_in(isec*NFIBERS+ifib).phi > 0 then
                            link_prev := '0';
                            link_next := '1';
                        elsif links_in(isec*NFIBERS+ifib).phi < 0 then
                            link_prev := '1';
                            link_next := '0';
                        else
                            link_prev := '0';
                            link_next := '0';
                        end if;
                    end if;
                    fifo_in(isec     *NFIFOS+ifib  ) <= links_in(isec*NFIBERS+ifib);
                    fifo_in(isec_next*NFIFOS+ifib+2).pt   <= links_in(isec*NFIBERS+ifib).pt;
                    fifo_in(isec_next*NFIFOS+ifib+2).eta  <= links_in(isec*NFIBERS+ifib).eta;
                    fifo_in(isec_next*NFIFOS+ifib+2).phi  <= links_in(isec*NFIBERS+ifib).phi - PHI_SHIFT;
                    fifo_in(isec_next*NFIFOS+ifib+2).rest <= links_in(isec*NFIBERS+ifib).rest;
                    fifo_in(isec_prev*NFIFOS+ifib+4).pt   <= links_in(isec*NFIBERS+ifib).pt;
                    fifo_in(isec_prev*NFIFOS+ifib+4).eta  <= links_in(isec*NFIBERS+ifib).eta;
                    fifo_in(isec_prev*NFIFOS+ifib+4).phi  <= links_in(isec*NFIBERS+ifib).phi + PHI_SHIFT;
                    fifo_in(isec_prev*NFIFOS+ifib+4).rest <= links_in(isec*NFIBERS+ifib).rest;
                    fifo_in_write(isec     *NFIFOS+ifib  ) <= link_this;
                    fifo_in_write(isec_next*NFIFOS+ifib+2) <= link_next;
                    fifo_in_write(isec_prev*NFIFOS+ifib+4) <= link_prev;
                    fifo_in_roll(isec     *NFIFOS+ifib  ) <= newevent;
                    fifo_in_roll(isec_next*NFIFOS+ifib+2) <= newevent;
                    fifo_in_roll(isec_prev*NFIFOS+ifib+4) <= newevent;
                end loop;
            end loop;
        end if;
    end process link2fifo;

    fifo2regions : process(ap_clk)
    begin
        if rising_edge(ap_clk) then
            for ireg in 0 to NREGIONS-1 loop
                if fifo_out_valid(ireg) = '1' then
                    regions_out(ireg) <= fifo_out(ireg);
                    regions_out_valid(ireg) <= '1';
                else
                    regions_out(ireg).pt   <= (others => '0');
                    regions_out(ireg).eta  <= (others => '0');
                    regions_out(ireg).phi  <= (others => '0');
                    regions_out(ireg).rest <= (others => '0');
                    regions_out_valid(ireg) <= '1';
                end if;
                regions_out_roll(ireg) <= fifo_out_roll(ireg);
            end loop;
        end if;
    end process fifo2regions;

    tracks_out_0_pt_V <= std_logic_vector(regions_out(0).pt);
    tracks_out_0_pt_V_ap_vld <= regions_out_valid(0);
    tracks_out_0_eta_V <= std_logic_vector(regions_out(0).eta);
    tracks_out_0_eta_V_ap_vld <= regions_out_valid(0);
    tracks_out_0_phi_V <= std_logic_vector(regions_out(0).phi);
    tracks_out_0_phi_V_ap_vld <= regions_out_valid(0);
    tracks_out_0_rest_V <= std_logic_vector(regions_out(0).rest);
    tracks_out_0_rest_V_ap_vld <= regions_out_valid(0);
    tracks_out_1_pt_V <= std_logic_vector(regions_out(1).pt);
    tracks_out_1_pt_V_ap_vld <= regions_out_valid(1);
    tracks_out_1_eta_V <= std_logic_vector(regions_out(1).eta);
    tracks_out_1_eta_V_ap_vld <= regions_out_valid(1);
    tracks_out_1_phi_V <= std_logic_vector(regions_out(1).phi);
    tracks_out_1_phi_V_ap_vld <= regions_out_valid(1);
    tracks_out_1_rest_V <= std_logic_vector(regions_out(1).rest);
    tracks_out_1_rest_V_ap_vld <= regions_out_valid(1);
    tracks_out_2_pt_V <= std_logic_vector(regions_out(2).pt);
    tracks_out_2_pt_V_ap_vld <= regions_out_valid(2);
    tracks_out_2_eta_V <= std_logic_vector(regions_out(2).eta);
    tracks_out_2_eta_V_ap_vld <= regions_out_valid(2);
    tracks_out_2_phi_V <= std_logic_vector(regions_out(2).phi);
    tracks_out_2_phi_V_ap_vld <= regions_out_valid(2);
    tracks_out_2_rest_V <= std_logic_vector(regions_out(2).rest);
    tracks_out_2_rest_V_ap_vld <= regions_out_valid(2);
    tracks_out_3_pt_V <= std_logic_vector(regions_out(3).pt);
    tracks_out_3_pt_V_ap_vld <= regions_out_valid(3);
    tracks_out_3_eta_V <= std_logic_vector(regions_out(3).eta);
    tracks_out_3_eta_V_ap_vld <= regions_out_valid(3);
    tracks_out_3_phi_V <= std_logic_vector(regions_out(3).phi);
    tracks_out_3_phi_V_ap_vld <= regions_out_valid(3);
    tracks_out_3_rest_V <= std_logic_vector(regions_out(3).rest);
    tracks_out_3_rest_V_ap_vld <= regions_out_valid(3);
    tracks_out_4_pt_V <= std_logic_vector(regions_out(4).pt);
    tracks_out_4_pt_V_ap_vld <= regions_out_valid(4);
    tracks_out_4_eta_V <= std_logic_vector(regions_out(4).eta);
    tracks_out_4_eta_V_ap_vld <= regions_out_valid(4);
    tracks_out_4_phi_V <= std_logic_vector(regions_out(4).phi);
    tracks_out_4_phi_V_ap_vld <= regions_out_valid(4);
    tracks_out_4_rest_V <= std_logic_vector(regions_out(4).rest);
    tracks_out_4_rest_V_ap_vld <= regions_out_valid(4);
    tracks_out_5_pt_V <= std_logic_vector(regions_out(5).pt);
    tracks_out_5_pt_V_ap_vld <= regions_out_valid(5);
    tracks_out_5_eta_V <= std_logic_vector(regions_out(5).eta);
    tracks_out_5_eta_V_ap_vld <= regions_out_valid(5);
    tracks_out_5_phi_V <= std_logic_vector(regions_out(5).phi);
    tracks_out_5_phi_V_ap_vld <= regions_out_valid(5);
    tracks_out_5_rest_V <= std_logic_vector(regions_out(5).rest);
    tracks_out_5_rest_V_ap_vld <= regions_out_valid(5);
    tracks_out_6_pt_V <= std_logic_vector(regions_out(6).pt);
    tracks_out_6_pt_V_ap_vld <= regions_out_valid(6);
    tracks_out_6_eta_V <= std_logic_vector(regions_out(6).eta);
    tracks_out_6_eta_V_ap_vld <= regions_out_valid(6);
    tracks_out_6_phi_V <= std_logic_vector(regions_out(6).phi);
    tracks_out_6_phi_V_ap_vld <= regions_out_valid(6);
    tracks_out_6_rest_V <= std_logic_vector(regions_out(6).rest);
    tracks_out_6_rest_V_ap_vld <= regions_out_valid(6);
    tracks_out_7_pt_V <= std_logic_vector(regions_out(7).pt);
    tracks_out_7_pt_V_ap_vld <= regions_out_valid(7);
    tracks_out_7_eta_V <= std_logic_vector(regions_out(7).eta);
    tracks_out_7_eta_V_ap_vld <= regions_out_valid(7);
    tracks_out_7_phi_V <= std_logic_vector(regions_out(7).phi);
    tracks_out_7_phi_V_ap_vld <= regions_out_valid(7);
    tracks_out_7_rest_V <= std_logic_vector(regions_out(7).rest);
    tracks_out_7_rest_V_ap_vld <= regions_out_valid(7);
    tracks_out_8_pt_V <= std_logic_vector(regions_out(8).pt);
    tracks_out_8_pt_V_ap_vld <= regions_out_valid(8);
    tracks_out_8_eta_V <= std_logic_vector(regions_out(8).eta);
    tracks_out_8_eta_V_ap_vld <= regions_out_valid(8);
    tracks_out_8_phi_V <= std_logic_vector(regions_out(8).phi);
    tracks_out_8_phi_V_ap_vld <= regions_out_valid(8);
    tracks_out_8_rest_V <= std_logic_vector(regions_out(8).rest);
    tracks_out_8_rest_V_ap_vld <= regions_out_valid(8);
    tracks_out_9_pt_V <= std_logic_vector(regions_out(9).pt);
    tracks_out_9_pt_V_ap_vld <= regions_out_valid(9);
    tracks_out_9_eta_V <= std_logic_vector(regions_out(9).eta);
    tracks_out_9_eta_V_ap_vld <= regions_out_valid(9);
    tracks_out_9_phi_V <= std_logic_vector(regions_out(9).phi);
    tracks_out_9_phi_V_ap_vld <= regions_out_valid(9);
    tracks_out_9_rest_V <= std_logic_vector(regions_out(9).rest);
    tracks_out_9_rest_V_ap_vld <= regions_out_valid(9);
    tracks_out_10_pt_V <= std_logic_vector(regions_out(10).pt);
    tracks_out_10_pt_V_ap_vld <= regions_out_valid(10);
    tracks_out_10_eta_V <= std_logic_vector(regions_out(10).eta);
    tracks_out_10_eta_V_ap_vld <= regions_out_valid(10);
    tracks_out_10_phi_V <= std_logic_vector(regions_out(10).phi);
    tracks_out_10_phi_V_ap_vld <= regions_out_valid(10);
    tracks_out_10_rest_V <= std_logic_vector(regions_out(10).rest);
    tracks_out_10_rest_V_ap_vld <= regions_out_valid(10);
    tracks_out_11_pt_V <= std_logic_vector(regions_out(11).pt);
    tracks_out_11_pt_V_ap_vld <= regions_out_valid(11);
    tracks_out_11_eta_V <= std_logic_vector(regions_out(11).eta);
    tracks_out_11_eta_V_ap_vld <= regions_out_valid(11);
    tracks_out_11_phi_V <= std_logic_vector(regions_out(11).phi);
    tracks_out_11_phi_V_ap_vld <= regions_out_valid(11);
    tracks_out_11_rest_V <= std_logic_vector(regions_out(11).rest);
    tracks_out_11_rest_V_ap_vld <= regions_out_valid(11);
    tracks_out_12_pt_V <= std_logic_vector(regions_out(12).pt);
    tracks_out_12_pt_V_ap_vld <= regions_out_valid(12);
    tracks_out_12_eta_V <= std_logic_vector(regions_out(12).eta);
    tracks_out_12_eta_V_ap_vld <= regions_out_valid(12);
    tracks_out_12_phi_V <= std_logic_vector(regions_out(12).phi);
    tracks_out_12_phi_V_ap_vld <= regions_out_valid(12);
    tracks_out_12_rest_V <= std_logic_vector(regions_out(12).rest);
    tracks_out_12_rest_V_ap_vld <= regions_out_valid(12);
    tracks_out_13_pt_V <= std_logic_vector(regions_out(13).pt);
    tracks_out_13_pt_V_ap_vld <= regions_out_valid(13);
    tracks_out_13_eta_V <= std_logic_vector(regions_out(13).eta);
    tracks_out_13_eta_V_ap_vld <= regions_out_valid(13);
    tracks_out_13_phi_V <= std_logic_vector(regions_out(13).phi);
    tracks_out_13_phi_V_ap_vld <= regions_out_valid(13);
    tracks_out_13_rest_V <= std_logic_vector(regions_out(13).rest);
    tracks_out_13_rest_V_ap_vld <= regions_out_valid(13);
    tracks_out_14_pt_V <= std_logic_vector(regions_out(14).pt);
    tracks_out_14_pt_V_ap_vld <= regions_out_valid(14);
    tracks_out_14_eta_V <= std_logic_vector(regions_out(14).eta);
    tracks_out_14_eta_V_ap_vld <= regions_out_valid(14);
    tracks_out_14_phi_V <= std_logic_vector(regions_out(14).phi);
    tracks_out_14_phi_V_ap_vld <= regions_out_valid(14);
    tracks_out_14_rest_V <= std_logic_vector(regions_out(14).rest);
    tracks_out_14_rest_V_ap_vld <= regions_out_valid(14);
    tracks_out_15_pt_V <= std_logic_vector(regions_out(15).pt);
    tracks_out_15_pt_V_ap_vld <= regions_out_valid(15);
    tracks_out_15_eta_V <= std_logic_vector(regions_out(15).eta);
    tracks_out_15_eta_V_ap_vld <= regions_out_valid(15);
    tracks_out_15_phi_V <= std_logic_vector(regions_out(15).phi);
    tracks_out_15_phi_V_ap_vld <= regions_out_valid(15);
    tracks_out_15_rest_V <= std_logic_vector(regions_out(15).rest);
    tracks_out_15_rest_V_ap_vld <= regions_out_valid(15);
    tracks_out_16_pt_V <= std_logic_vector(regions_out(16).pt);
    tracks_out_16_pt_V_ap_vld <= regions_out_valid(16);
    tracks_out_16_eta_V <= std_logic_vector(regions_out(16).eta);
    tracks_out_16_eta_V_ap_vld <= regions_out_valid(16);
    tracks_out_16_phi_V <= std_logic_vector(regions_out(16).phi);
    tracks_out_16_phi_V_ap_vld <= regions_out_valid(16);
    tracks_out_16_rest_V <= std_logic_vector(regions_out(16).rest);
    tracks_out_16_rest_V_ap_vld <= regions_out_valid(16);
    tracks_out_17_pt_V <= std_logic_vector(regions_out(17).pt);
    tracks_out_17_pt_V_ap_vld <= regions_out_valid(17);
    tracks_out_17_eta_V <= std_logic_vector(regions_out(17).eta);
    tracks_out_17_eta_V_ap_vld <= regions_out_valid(17);
    tracks_out_17_phi_V <= std_logic_vector(regions_out(17).phi);
    tracks_out_17_phi_V_ap_vld <= regions_out_valid(17);
    tracks_out_17_rest_V <= std_logic_vector(regions_out(17).rest);
    tracks_out_17_rest_V_ap_vld <= regions_out_valid(17);
    tracks_out_18_pt_V <= std_logic_vector(regions_out(18).pt);
    tracks_out_18_pt_V_ap_vld <= regions_out_valid(18);
    tracks_out_18_eta_V <= std_logic_vector(regions_out(18).eta);
    tracks_out_18_eta_V_ap_vld <= regions_out_valid(18);
    tracks_out_18_phi_V <= std_logic_vector(regions_out(18).phi);
    tracks_out_18_phi_V_ap_vld <= regions_out_valid(18);
    tracks_out_18_rest_V <= std_logic_vector(regions_out(18).rest);
    tracks_out_18_rest_V_ap_vld <= regions_out_valid(18);
    tracks_out_19_pt_V <= std_logic_vector(regions_out(19).pt);
    tracks_out_19_pt_V_ap_vld <= regions_out_valid(19);
    tracks_out_19_eta_V <= std_logic_vector(regions_out(19).eta);
    tracks_out_19_eta_V_ap_vld <= regions_out_valid(19);
    tracks_out_19_phi_V <= std_logic_vector(regions_out(19).phi);
    tracks_out_19_phi_V_ap_vld <= regions_out_valid(19);
    tracks_out_19_rest_V <= std_logic_vector(regions_out(19).rest);
    tracks_out_19_rest_V_ap_vld <= regions_out_valid(19);
    tracks_out_20_pt_V <= std_logic_vector(regions_out(20).pt);
    tracks_out_20_pt_V_ap_vld <= regions_out_valid(20);
    tracks_out_20_eta_V <= std_logic_vector(regions_out(20).eta);
    tracks_out_20_eta_V_ap_vld <= regions_out_valid(20);
    tracks_out_20_phi_V <= std_logic_vector(regions_out(20).phi);
    tracks_out_20_phi_V_ap_vld <= regions_out_valid(20);
    tracks_out_20_rest_V <= std_logic_vector(regions_out(20).rest);
    tracks_out_20_rest_V_ap_vld <= regions_out_valid(20);
    tracks_out_21_pt_V <= std_logic_vector(regions_out(21).pt);
    tracks_out_21_pt_V_ap_vld <= regions_out_valid(21);
    tracks_out_21_eta_V <= std_logic_vector(regions_out(21).eta);
    tracks_out_21_eta_V_ap_vld <= regions_out_valid(21);
    tracks_out_21_phi_V <= std_logic_vector(regions_out(21).phi);
    tracks_out_21_phi_V_ap_vld <= regions_out_valid(21);
    tracks_out_21_rest_V <= std_logic_vector(regions_out(21).rest);
    tracks_out_21_rest_V_ap_vld <= regions_out_valid(21);
    tracks_out_22_pt_V <= std_logic_vector(regions_out(22).pt);
    tracks_out_22_pt_V_ap_vld <= regions_out_valid(22);
    tracks_out_22_eta_V <= std_logic_vector(regions_out(22).eta);
    tracks_out_22_eta_V_ap_vld <= regions_out_valid(22);
    tracks_out_22_phi_V <= std_logic_vector(regions_out(22).phi);
    tracks_out_22_phi_V_ap_vld <= regions_out_valid(22);
    tracks_out_22_rest_V <= std_logic_vector(regions_out(22).rest);
    tracks_out_22_rest_V_ap_vld <= regions_out_valid(22);
    tracks_out_23_pt_V <= std_logic_vector(regions_out(23).pt);
    tracks_out_23_pt_V_ap_vld <= regions_out_valid(23);
    tracks_out_23_eta_V <= std_logic_vector(regions_out(23).eta);
    tracks_out_23_eta_V_ap_vld <= regions_out_valid(23);
    tracks_out_23_phi_V <= std_logic_vector(regions_out(23).phi);
    tracks_out_23_phi_V_ap_vld <= regions_out_valid(23);
    tracks_out_23_rest_V <= std_logic_vector(regions_out(23).rest);
    tracks_out_23_rest_V_ap_vld <= regions_out_valid(23);
    tracks_out_24_pt_V <= std_logic_vector(regions_out(24).pt);
    tracks_out_24_pt_V_ap_vld <= regions_out_valid(24);
    tracks_out_24_eta_V <= std_logic_vector(regions_out(24).eta);
    tracks_out_24_eta_V_ap_vld <= regions_out_valid(24);
    tracks_out_24_phi_V <= std_logic_vector(regions_out(24).phi);
    tracks_out_24_phi_V_ap_vld <= regions_out_valid(24);
    tracks_out_24_rest_V <= std_logic_vector(regions_out(24).rest);
    tracks_out_24_rest_V_ap_vld <= regions_out_valid(24);
    tracks_out_25_pt_V <= std_logic_vector(regions_out(25).pt);
    tracks_out_25_pt_V_ap_vld <= regions_out_valid(25);
    tracks_out_25_eta_V <= std_logic_vector(regions_out(25).eta);
    tracks_out_25_eta_V_ap_vld <= regions_out_valid(25);
    tracks_out_25_phi_V <= std_logic_vector(regions_out(25).phi);
    tracks_out_25_phi_V_ap_vld <= regions_out_valid(25);
    tracks_out_25_rest_V <= std_logic_vector(regions_out(25).rest);
    tracks_out_25_rest_V_ap_vld <= regions_out_valid(25);
    tracks_out_26_pt_V <= std_logic_vector(regions_out(26).pt);
    tracks_out_26_pt_V_ap_vld <= regions_out_valid(26);
    tracks_out_26_eta_V <= std_logic_vector(regions_out(26).eta);
    tracks_out_26_eta_V_ap_vld <= regions_out_valid(26);
    tracks_out_26_phi_V <= std_logic_vector(regions_out(26).phi);
    tracks_out_26_phi_V_ap_vld <= regions_out_valid(26);
    tracks_out_26_rest_V <= std_logic_vector(regions_out(26).rest);
    tracks_out_26_rest_V_ap_vld <= regions_out_valid(26);
    tracks_out_27_pt_V <= std_logic_vector(regions_out(27).pt);
    tracks_out_27_pt_V_ap_vld <= regions_out_valid(27);
    tracks_out_27_eta_V <= std_logic_vector(regions_out(27).eta);
    tracks_out_27_eta_V_ap_vld <= regions_out_valid(27);
    tracks_out_27_phi_V <= std_logic_vector(regions_out(27).phi);
    tracks_out_27_phi_V_ap_vld <= regions_out_valid(27);
    tracks_out_27_rest_V <= std_logic_vector(regions_out(27).rest);
    tracks_out_27_rest_V_ap_vld <= regions_out_valid(27);
    tracks_out_28_pt_V <= std_logic_vector(regions_out(28).pt);
    tracks_out_28_pt_V_ap_vld <= regions_out_valid(28);
    tracks_out_28_eta_V <= std_logic_vector(regions_out(28).eta);
    tracks_out_28_eta_V_ap_vld <= regions_out_valid(28);
    tracks_out_28_phi_V <= std_logic_vector(regions_out(28).phi);
    tracks_out_28_phi_V_ap_vld <= regions_out_valid(28);
    tracks_out_28_rest_V <= std_logic_vector(regions_out(28).rest);
    tracks_out_28_rest_V_ap_vld <= regions_out_valid(28);
    tracks_out_29_pt_V <= std_logic_vector(regions_out(29).pt);
    tracks_out_29_pt_V_ap_vld <= regions_out_valid(29);
    tracks_out_29_eta_V <= std_logic_vector(regions_out(29).eta);
    tracks_out_29_eta_V_ap_vld <= regions_out_valid(29);
    tracks_out_29_phi_V <= std_logic_vector(regions_out(29).phi);
    tracks_out_29_phi_V_ap_vld <= regions_out_valid(29);
    tracks_out_29_rest_V <= std_logic_vector(regions_out(29).rest);
    tracks_out_29_rest_V_ap_vld <= regions_out_valid(29);
    tracks_out_30_pt_V <= std_logic_vector(regions_out(30).pt);
    tracks_out_30_pt_V_ap_vld <= regions_out_valid(30);
    tracks_out_30_eta_V <= std_logic_vector(regions_out(30).eta);
    tracks_out_30_eta_V_ap_vld <= regions_out_valid(30);
    tracks_out_30_phi_V <= std_logic_vector(regions_out(30).phi);
    tracks_out_30_phi_V_ap_vld <= regions_out_valid(30);
    tracks_out_30_rest_V <= std_logic_vector(regions_out(30).rest);
    tracks_out_30_rest_V_ap_vld <= regions_out_valid(30);
    tracks_out_31_pt_V <= std_logic_vector(regions_out(31).pt);
    tracks_out_31_pt_V_ap_vld <= regions_out_valid(31);
    tracks_out_31_eta_V <= std_logic_vector(regions_out(31).eta);
    tracks_out_31_eta_V_ap_vld <= regions_out_valid(31);
    tracks_out_31_phi_V <= std_logic_vector(regions_out(31).phi);
    tracks_out_31_phi_V_ap_vld <= regions_out_valid(31);
    tracks_out_31_rest_V <= std_logic_vector(regions_out(31).rest);
    tracks_out_31_rest_V_ap_vld <= regions_out_valid(31);
    tracks_out_32_pt_V <= std_logic_vector(regions_out(32).pt);
    tracks_out_32_pt_V_ap_vld <= regions_out_valid(32);
    tracks_out_32_eta_V <= std_logic_vector(regions_out(32).eta);
    tracks_out_32_eta_V_ap_vld <= regions_out_valid(32);
    tracks_out_32_phi_V <= std_logic_vector(regions_out(32).phi);
    tracks_out_32_phi_V_ap_vld <= regions_out_valid(32);
    tracks_out_32_rest_V <= std_logic_vector(regions_out(32).rest);
    tracks_out_32_rest_V_ap_vld <= regions_out_valid(32);
    tracks_out_33_pt_V <= std_logic_vector(regions_out(33).pt);
    tracks_out_33_pt_V_ap_vld <= regions_out_valid(33);
    tracks_out_33_eta_V <= std_logic_vector(regions_out(33).eta);
    tracks_out_33_eta_V_ap_vld <= regions_out_valid(33);
    tracks_out_33_phi_V <= std_logic_vector(regions_out(33).phi);
    tracks_out_33_phi_V_ap_vld <= regions_out_valid(33);
    tracks_out_33_rest_V <= std_logic_vector(regions_out(33).rest);
    tracks_out_33_rest_V_ap_vld <= regions_out_valid(33);
    tracks_out_34_pt_V <= std_logic_vector(regions_out(34).pt);
    tracks_out_34_pt_V_ap_vld <= regions_out_valid(34);
    tracks_out_34_eta_V <= std_logic_vector(regions_out(34).eta);
    tracks_out_34_eta_V_ap_vld <= regions_out_valid(34);
    tracks_out_34_phi_V <= std_logic_vector(regions_out(34).phi);
    tracks_out_34_phi_V_ap_vld <= regions_out_valid(34);
    tracks_out_34_rest_V <= std_logic_vector(regions_out(34).rest);
    tracks_out_34_rest_V_ap_vld <= regions_out_valid(34);
    tracks_out_35_pt_V <= std_logic_vector(regions_out(35).pt);
    tracks_out_35_pt_V_ap_vld <= regions_out_valid(35);
    tracks_out_35_eta_V <= std_logic_vector(regions_out(35).eta);
    tracks_out_35_eta_V_ap_vld <= regions_out_valid(35);
    tracks_out_35_phi_V <= std_logic_vector(regions_out(35).phi);
    tracks_out_35_phi_V_ap_vld <= regions_out_valid(35);
    tracks_out_35_rest_V <= std_logic_vector(regions_out(35).rest);
    tracks_out_35_rest_V_ap_vld <= regions_out_valid(35);
    tracks_out_36_pt_V <= std_logic_vector(regions_out(36).pt);
    tracks_out_36_pt_V_ap_vld <= regions_out_valid(36);
    tracks_out_36_eta_V <= std_logic_vector(regions_out(36).eta);
    tracks_out_36_eta_V_ap_vld <= regions_out_valid(36);
    tracks_out_36_phi_V <= std_logic_vector(regions_out(36).phi);
    tracks_out_36_phi_V_ap_vld <= regions_out_valid(36);
    tracks_out_36_rest_V <= std_logic_vector(regions_out(36).rest);
    tracks_out_36_rest_V_ap_vld <= regions_out_valid(36);
    tracks_out_37_pt_V <= std_logic_vector(regions_out(37).pt);
    tracks_out_37_pt_V_ap_vld <= regions_out_valid(37);
    tracks_out_37_eta_V <= std_logic_vector(regions_out(37).eta);
    tracks_out_37_eta_V_ap_vld <= regions_out_valid(37);
    tracks_out_37_phi_V <= std_logic_vector(regions_out(37).phi);
    tracks_out_37_phi_V_ap_vld <= regions_out_valid(37);
    tracks_out_37_rest_V <= std_logic_vector(regions_out(37).rest);
    tracks_out_37_rest_V_ap_vld <= regions_out_valid(37);
    tracks_out_38_pt_V <= std_logic_vector(regions_out(38).pt);
    tracks_out_38_pt_V_ap_vld <= regions_out_valid(38);
    tracks_out_38_eta_V <= std_logic_vector(regions_out(38).eta);
    tracks_out_38_eta_V_ap_vld <= regions_out_valid(38);
    tracks_out_38_phi_V <= std_logic_vector(regions_out(38).phi);
    tracks_out_38_phi_V_ap_vld <= regions_out_valid(38);
    tracks_out_38_rest_V <= std_logic_vector(regions_out(38).rest);
    tracks_out_38_rest_V_ap_vld <= regions_out_valid(38);
    tracks_out_39_pt_V <= std_logic_vector(regions_out(39).pt);
    tracks_out_39_pt_V_ap_vld <= regions_out_valid(39);
    tracks_out_39_eta_V <= std_logic_vector(regions_out(39).eta);
    tracks_out_39_eta_V_ap_vld <= regions_out_valid(39);
    tracks_out_39_phi_V <= std_logic_vector(regions_out(39).phi);
    tracks_out_39_phi_V_ap_vld <= regions_out_valid(39);
    tracks_out_39_rest_V <= std_logic_vector(regions_out(39).rest);
    tracks_out_39_rest_V_ap_vld <= regions_out_valid(39);
    tracks_out_40_pt_V <= std_logic_vector(regions_out(40).pt);
    tracks_out_40_pt_V_ap_vld <= regions_out_valid(40);
    tracks_out_40_eta_V <= std_logic_vector(regions_out(40).eta);
    tracks_out_40_eta_V_ap_vld <= regions_out_valid(40);
    tracks_out_40_phi_V <= std_logic_vector(regions_out(40).phi);
    tracks_out_40_phi_V_ap_vld <= regions_out_valid(40);
    tracks_out_40_rest_V <= std_logic_vector(regions_out(40).rest);
    tracks_out_40_rest_V_ap_vld <= regions_out_valid(40);
    tracks_out_41_pt_V <= std_logic_vector(regions_out(41).pt);
    tracks_out_41_pt_V_ap_vld <= regions_out_valid(41);
    tracks_out_41_eta_V <= std_logic_vector(regions_out(41).eta);
    tracks_out_41_eta_V_ap_vld <= regions_out_valid(41);
    tracks_out_41_phi_V <= std_logic_vector(regions_out(41).phi);
    tracks_out_41_phi_V_ap_vld <= regions_out_valid(41);
    tracks_out_41_rest_V <= std_logic_vector(regions_out(41).rest);
    tracks_out_41_rest_V_ap_vld <= regions_out_valid(41);
    tracks_out_42_pt_V <= std_logic_vector(regions_out(42).pt);
    tracks_out_42_pt_V_ap_vld <= regions_out_valid(42);
    tracks_out_42_eta_V <= std_logic_vector(regions_out(42).eta);
    tracks_out_42_eta_V_ap_vld <= regions_out_valid(42);
    tracks_out_42_phi_V <= std_logic_vector(regions_out(42).phi);
    tracks_out_42_phi_V_ap_vld <= regions_out_valid(42);
    tracks_out_42_rest_V <= std_logic_vector(regions_out(42).rest);
    tracks_out_42_rest_V_ap_vld <= regions_out_valid(42);
    tracks_out_43_pt_V <= std_logic_vector(regions_out(43).pt);
    tracks_out_43_pt_V_ap_vld <= regions_out_valid(43);
    tracks_out_43_eta_V <= std_logic_vector(regions_out(43).eta);
    tracks_out_43_eta_V_ap_vld <= regions_out_valid(43);
    tracks_out_43_phi_V <= std_logic_vector(regions_out(43).phi);
    tracks_out_43_phi_V_ap_vld <= regions_out_valid(43);
    tracks_out_43_rest_V <= std_logic_vector(regions_out(43).rest);
    tracks_out_43_rest_V_ap_vld <= regions_out_valid(43);
    tracks_out_44_pt_V <= std_logic_vector(regions_out(44).pt);
    tracks_out_44_pt_V_ap_vld <= regions_out_valid(44);
    tracks_out_44_eta_V <= std_logic_vector(regions_out(44).eta);
    tracks_out_44_eta_V_ap_vld <= regions_out_valid(44);
    tracks_out_44_phi_V <= std_logic_vector(regions_out(44).phi);
    tracks_out_44_phi_V_ap_vld <= regions_out_valid(44);
    tracks_out_44_rest_V <= std_logic_vector(regions_out(44).rest);
    tracks_out_44_rest_V_ap_vld <= regions_out_valid(44);
    tracks_out_45_pt_V <= std_logic_vector(regions_out(45).pt);
    tracks_out_45_pt_V_ap_vld <= regions_out_valid(45);
    tracks_out_45_eta_V <= std_logic_vector(regions_out(45).eta);
    tracks_out_45_eta_V_ap_vld <= regions_out_valid(45);
    tracks_out_45_phi_V <= std_logic_vector(regions_out(45).phi);
    tracks_out_45_phi_V_ap_vld <= regions_out_valid(45);
    tracks_out_45_rest_V <= std_logic_vector(regions_out(45).rest);
    tracks_out_45_rest_V_ap_vld <= regions_out_valid(45);
    tracks_out_46_pt_V <= std_logic_vector(regions_out(46).pt);
    tracks_out_46_pt_V_ap_vld <= regions_out_valid(46);
    tracks_out_46_eta_V <= std_logic_vector(regions_out(46).eta);
    tracks_out_46_eta_V_ap_vld <= regions_out_valid(46);
    tracks_out_46_phi_V <= std_logic_vector(regions_out(46).phi);
    tracks_out_46_phi_V_ap_vld <= regions_out_valid(46);
    tracks_out_46_rest_V <= std_logic_vector(regions_out(46).rest);
    tracks_out_46_rest_V_ap_vld <= regions_out_valid(46);
    tracks_out_47_pt_V <= std_logic_vector(regions_out(47).pt);
    tracks_out_47_pt_V_ap_vld <= regions_out_valid(47);
    tracks_out_47_eta_V <= std_logic_vector(regions_out(47).eta);
    tracks_out_47_eta_V_ap_vld <= regions_out_valid(47);
    tracks_out_47_phi_V <= std_logic_vector(regions_out(47).phi);
    tracks_out_47_phi_V_ap_vld <= regions_out_valid(47);
    tracks_out_47_rest_V <= std_logic_vector(regions_out(47).rest);
    tracks_out_47_rest_V_ap_vld <= regions_out_valid(47);
    tracks_out_48_pt_V <= std_logic_vector(regions_out(48).pt);
    tracks_out_48_pt_V_ap_vld <= regions_out_valid(48);
    tracks_out_48_eta_V <= std_logic_vector(regions_out(48).eta);
    tracks_out_48_eta_V_ap_vld <= regions_out_valid(48);
    tracks_out_48_phi_V <= std_logic_vector(regions_out(48).phi);
    tracks_out_48_phi_V_ap_vld <= regions_out_valid(48);
    tracks_out_48_rest_V <= std_logic_vector(regions_out(48).rest);
    tracks_out_48_rest_V_ap_vld <= regions_out_valid(48);
    tracks_out_49_pt_V <= std_logic_vector(regions_out(49).pt);
    tracks_out_49_pt_V_ap_vld <= regions_out_valid(49);
    tracks_out_49_eta_V <= std_logic_vector(regions_out(49).eta);
    tracks_out_49_eta_V_ap_vld <= regions_out_valid(49);
    tracks_out_49_phi_V <= std_logic_vector(regions_out(49).phi);
    tracks_out_49_phi_V_ap_vld <= regions_out_valid(49);
    tracks_out_49_rest_V <= std_logic_vector(regions_out(49).rest);
    tracks_out_49_rest_V_ap_vld <= regions_out_valid(49);
    tracks_out_50_pt_V <= std_logic_vector(regions_out(50).pt);
    tracks_out_50_pt_V_ap_vld <= regions_out_valid(50);
    tracks_out_50_eta_V <= std_logic_vector(regions_out(50).eta);
    tracks_out_50_eta_V_ap_vld <= regions_out_valid(50);
    tracks_out_50_phi_V <= std_logic_vector(regions_out(50).phi);
    tracks_out_50_phi_V_ap_vld <= regions_out_valid(50);
    tracks_out_50_rest_V <= std_logic_vector(regions_out(50).rest);
    tracks_out_50_rest_V_ap_vld <= regions_out_valid(50);
    tracks_out_51_pt_V <= std_logic_vector(regions_out(51).pt);
    tracks_out_51_pt_V_ap_vld <= regions_out_valid(51);
    tracks_out_51_eta_V <= std_logic_vector(regions_out(51).eta);
    tracks_out_51_eta_V_ap_vld <= regions_out_valid(51);
    tracks_out_51_phi_V <= std_logic_vector(regions_out(51).phi);
    tracks_out_51_phi_V_ap_vld <= regions_out_valid(51);
    tracks_out_51_rest_V <= std_logic_vector(regions_out(51).rest);
    tracks_out_51_rest_V_ap_vld <= regions_out_valid(51);
    tracks_out_52_pt_V <= std_logic_vector(regions_out(52).pt);
    tracks_out_52_pt_V_ap_vld <= regions_out_valid(52);
    tracks_out_52_eta_V <= std_logic_vector(regions_out(52).eta);
    tracks_out_52_eta_V_ap_vld <= regions_out_valid(52);
    tracks_out_52_phi_V <= std_logic_vector(regions_out(52).phi);
    tracks_out_52_phi_V_ap_vld <= regions_out_valid(52);
    tracks_out_52_rest_V <= std_logic_vector(regions_out(52).rest);
    tracks_out_52_rest_V_ap_vld <= regions_out_valid(52);
    tracks_out_53_pt_V <= std_logic_vector(regions_out(53).pt);
    tracks_out_53_pt_V_ap_vld <= regions_out_valid(53);
    tracks_out_53_eta_V <= std_logic_vector(regions_out(53).eta);
    tracks_out_53_eta_V_ap_vld <= regions_out_valid(53);
    tracks_out_53_phi_V <= std_logic_vector(regions_out(53).phi);
    tracks_out_53_phi_V_ap_vld <= regions_out_valid(53);
    tracks_out_53_rest_V <= std_logic_vector(regions_out(53).rest);
    tracks_out_53_rest_V_ap_vld <= regions_out_valid(53);
    newevent_out <= regions_out_roll(0);

end Behavioral;
