library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.regionizer_data.all;

entity calo_regionizer is
    port(
            ap_clk : IN STD_LOGIC;
            ap_rst : IN STD_LOGIC;
            ap_start : IN STD_LOGIC;
            ap_done : OUT STD_LOGIC;
            ap_idle : OUT STD_LOGIC;
            ap_ready : OUT STD_LOGIC;
            newevent : IN STD_LOGIC;
            tracks_in_0_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_0_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_0_2_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_2_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_2_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_2_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_0_3_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_3_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_3_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_3_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_2_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_2_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_2_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_2_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_3_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_3_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_3_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_3_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_2_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_2_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_2_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_2_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_3_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_3_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_3_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_3_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_0_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_0_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_1_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_1_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_2_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_2_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_3_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_3_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_4_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_4_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_5_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_5_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_6_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_6_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_7_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_7_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_8_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_8_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            newevent_out : OUT STD_LOGIC

    );
end calo_regionizer;

architecture Behavioral of calo_regionizer is
    constant NREGIONS  : natural := NSECTORS;
    constant NALLFIFOS : natural := NCALOSECTORS*NCALOFIFOS;
    constant NMERGE2   : natural := NALLFIFOS/2;
    constant NMERGE4   : natural := NALLFIFOS/4;

    signal links_in :       particles(NCALOSECTORS*NCALOFIBERS-1 downto 0);
    signal fifo_in :        particles(NALLFIFOS-1 downto 0);
    signal fifo_write :     std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');

    signal fifo_out :         particles(NALLFIFOS-1 downto 0);
    signal fifo_out_valid :   std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');
    signal fifo_full:         std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');
    signal fifo_out_roll:     std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');

    signal merged2_out :        particles(NMERGE2-1 downto 0);
    signal merged2_out_valid :  std_logic_vector(NMERGE2-1 downto 0) := (others => '0');
    signal merged2_out_roll:    std_logic_vector(NMERGE2-1 downto 0) := (others => '0');
    signal merged2_full:        std_logic_vector(NMERGE2-1 downto 0) := (others => '0');

    signal merged4_out :        particles(NMERGE4-1 downto 0);
    signal merged4_out_valid :  std_logic_vector(NMERGE4-1 downto 0) := (others => '0');
    signal merged4_out_roll:    std_logic_vector(NMERGE4-1 downto 0) := (others => '0');
    signal merged4_full:        std_logic_vector(NMERGE4-1 downto 0) := (others => '0');

    signal merged_out :        particles(NREGIONS-1 downto 0);
    signal merged_out_valid :  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal merged_out_roll:    std_logic_vector(NREGIONS-1 downto 0) := (others => '0');

    signal newevent_del : std_logic;
begin

    delay : process (ap_clk)
    begin
        if rising_edge(ap_clk) then
            newevent_del <= newevent;
        end if;
    end process delay;

    input_slice : entity work.calo_router_input_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     tracks_in_0_0_eta_V => tracks_in_0_0_eta_V,
                     tracks_in_0_0_phi_V => tracks_in_0_0_phi_V,
                     tracks_in_0_0_pt_V => tracks_in_0_0_pt_V,
                     tracks_in_0_0_rest_V => tracks_in_0_0_rest_V,
                     tracks_in_0_1_eta_V => tracks_in_0_1_eta_V,
                     tracks_in_0_1_phi_V => tracks_in_0_1_phi_V,
                     tracks_in_0_1_pt_V => tracks_in_0_1_pt_V,
                     tracks_in_0_1_rest_V => tracks_in_0_1_rest_V,
                     tracks_in_0_2_eta_V => tracks_in_0_2_eta_V,
                     tracks_in_0_2_phi_V => tracks_in_0_2_phi_V,
                     tracks_in_0_2_pt_V => tracks_in_0_2_pt_V,
                     tracks_in_0_2_rest_V => tracks_in_0_2_rest_V,
                     tracks_in_0_3_eta_V => tracks_in_0_3_eta_V,
                     tracks_in_0_3_phi_V => tracks_in_0_3_phi_V,
                     tracks_in_0_3_pt_V => tracks_in_0_3_pt_V,
                     tracks_in_0_3_rest_V => tracks_in_0_3_rest_V,
                     tracks_in_1_0_eta_V => tracks_in_1_0_eta_V,
                     tracks_in_1_0_phi_V => tracks_in_1_0_phi_V,
                     tracks_in_1_0_pt_V => tracks_in_1_0_pt_V,
                     tracks_in_1_0_rest_V => tracks_in_1_0_rest_V,
                     tracks_in_1_1_eta_V => tracks_in_1_1_eta_V,
                     tracks_in_1_1_phi_V => tracks_in_1_1_phi_V,
                     tracks_in_1_1_pt_V => tracks_in_1_1_pt_V,
                     tracks_in_1_1_rest_V => tracks_in_1_1_rest_V,
                     tracks_in_1_2_eta_V => tracks_in_1_2_eta_V,
                     tracks_in_1_2_phi_V => tracks_in_1_2_phi_V,
                     tracks_in_1_2_pt_V => tracks_in_1_2_pt_V,
                     tracks_in_1_2_rest_V => tracks_in_1_2_rest_V,
                     tracks_in_1_3_eta_V => tracks_in_1_3_eta_V,
                     tracks_in_1_3_phi_V => tracks_in_1_3_phi_V,
                     tracks_in_1_3_pt_V => tracks_in_1_3_pt_V,
                     tracks_in_1_3_rest_V => tracks_in_1_3_rest_V,
                     tracks_in_2_0_eta_V => tracks_in_2_0_eta_V,
                     tracks_in_2_0_phi_V => tracks_in_2_0_phi_V,
                     tracks_in_2_0_pt_V => tracks_in_2_0_pt_V,
                     tracks_in_2_0_rest_V => tracks_in_2_0_rest_V,
                     tracks_in_2_1_eta_V => tracks_in_2_1_eta_V,
                     tracks_in_2_1_phi_V => tracks_in_2_1_phi_V,
                     tracks_in_2_1_pt_V => tracks_in_2_1_pt_V,
                     tracks_in_2_1_rest_V => tracks_in_2_1_rest_V,
                     tracks_in_2_2_eta_V => tracks_in_2_2_eta_V,
                     tracks_in_2_2_phi_V => tracks_in_2_2_phi_V,
                     tracks_in_2_2_pt_V => tracks_in_2_2_pt_V,
                     tracks_in_2_2_rest_V => tracks_in_2_2_rest_V,
                     tracks_in_2_3_eta_V => tracks_in_2_3_eta_V,
                     tracks_in_2_3_phi_V => tracks_in_2_3_phi_V,
                     tracks_in_2_3_pt_V => tracks_in_2_3_pt_V,
                     tracks_in_2_3_rest_V => tracks_in_2_3_rest_V,
                     fifo_in_0_0_pt_V  => fifo_in(0*NCALOFIFOS+ 0).pt,
                     fifo_in_0_1_pt_V  => fifo_in(0*NCALOFIFOS+ 1).pt,
                     fifo_in_0_2_pt_V  => fifo_in(0*NCALOFIFOS+ 2).pt,
                     fifo_in_0_3_pt_V  => fifo_in(0*NCALOFIFOS+ 3).pt,
                     fifo_in_0_4_pt_V  => fifo_in(0*NCALOFIFOS+ 4).pt,
                     fifo_in_0_5_pt_V  => fifo_in(0*NCALOFIFOS+ 5).pt,
                     fifo_in_0_6_pt_V  => fifo_in(0*NCALOFIFOS+ 6).pt,
                     fifo_in_0_7_pt_V  => fifo_in(0*NCALOFIFOS+ 7).pt,
                     fifo_in_0_8_pt_V  => fifo_in(0*NCALOFIFOS+ 8).pt,
                     fifo_in_0_9_pt_V  => fifo_in(0*NCALOFIFOS+ 9).pt,
                     fifo_in_0_10_pt_V => fifo_in(0*NCALOFIFOS+10).pt,
                     fifo_in_0_11_pt_V => fifo_in(0*NCALOFIFOS+11).pt,
                     fifo_in_0_12_pt_V => fifo_in(0*NCALOFIFOS+12).pt,
                     fifo_in_0_13_pt_V => fifo_in(0*NCALOFIFOS+13).pt,
                     fifo_in_0_14_pt_V => fifo_in(0*NCALOFIFOS+14).pt,
                     fifo_in_0_15_pt_V => fifo_in(0*NCALOFIFOS+15).pt,
                     fifo_in_0_16_pt_V => fifo_in(0*NCALOFIFOS+16).pt,
                     fifo_in_0_17_pt_V => fifo_in(0*NCALOFIFOS+17).pt,
                     fifo_in_0_18_pt_V => fifo_in(0*NCALOFIFOS+18).pt,
                     fifo_in_0_19_pt_V => fifo_in(0*NCALOFIFOS+19).pt,
                     fifo_in_1_0_pt_V  => fifo_in(1*NCALOFIFOS+ 0).pt,
                     fifo_in_1_1_pt_V  => fifo_in(1*NCALOFIFOS+ 1).pt,
                     fifo_in_1_2_pt_V  => fifo_in(1*NCALOFIFOS+ 2).pt,
                     fifo_in_1_3_pt_V  => fifo_in(1*NCALOFIFOS+ 3).pt,
                     fifo_in_1_4_pt_V  => fifo_in(1*NCALOFIFOS+ 4).pt,
                     fifo_in_1_5_pt_V  => fifo_in(1*NCALOFIFOS+ 5).pt,
                     fifo_in_1_6_pt_V  => fifo_in(1*NCALOFIFOS+ 6).pt,
                     fifo_in_1_7_pt_V  => fifo_in(1*NCALOFIFOS+ 7).pt,
                     fifo_in_1_8_pt_V  => fifo_in(1*NCALOFIFOS+ 8).pt,
                     fifo_in_1_9_pt_V  => fifo_in(1*NCALOFIFOS+ 9).pt,
                     fifo_in_1_10_pt_V => fifo_in(1*NCALOFIFOS+10).pt,
                     fifo_in_1_11_pt_V => fifo_in(1*NCALOFIFOS+11).pt,
                     fifo_in_1_12_pt_V => fifo_in(1*NCALOFIFOS+12).pt,
                     fifo_in_1_13_pt_V => fifo_in(1*NCALOFIFOS+13).pt,
                     fifo_in_1_14_pt_V => fifo_in(1*NCALOFIFOS+14).pt,
                     fifo_in_1_15_pt_V => fifo_in(1*NCALOFIFOS+15).pt,
                     fifo_in_1_16_pt_V => fifo_in(1*NCALOFIFOS+16).pt,
                     fifo_in_1_17_pt_V => fifo_in(1*NCALOFIFOS+17).pt,
                     fifo_in_1_18_pt_V => fifo_in(1*NCALOFIFOS+18).pt,
                     fifo_in_1_19_pt_V => fifo_in(1*NCALOFIFOS+19).pt,
                     fifo_in_2_0_pt_V  => fifo_in(2*NCALOFIFOS+ 0).pt,
                     fifo_in_2_1_pt_V  => fifo_in(2*NCALOFIFOS+ 1).pt,
                     fifo_in_2_2_pt_V  => fifo_in(2*NCALOFIFOS+ 2).pt,
                     fifo_in_2_3_pt_V  => fifo_in(2*NCALOFIFOS+ 3).pt,
                     fifo_in_2_4_pt_V  => fifo_in(2*NCALOFIFOS+ 4).pt,
                     fifo_in_2_5_pt_V  => fifo_in(2*NCALOFIFOS+ 5).pt,
                     fifo_in_2_6_pt_V  => fifo_in(2*NCALOFIFOS+ 6).pt,
                     fifo_in_2_7_pt_V  => fifo_in(2*NCALOFIFOS+ 7).pt,
                     fifo_in_2_8_pt_V  => fifo_in(2*NCALOFIFOS+ 8).pt,
                     fifo_in_2_9_pt_V  => fifo_in(2*NCALOFIFOS+ 9).pt,
                     fifo_in_2_10_pt_V => fifo_in(2*NCALOFIFOS+10).pt,
                     fifo_in_2_11_pt_V => fifo_in(2*NCALOFIFOS+11).pt,
                     fifo_in_2_12_pt_V => fifo_in(2*NCALOFIFOS+12).pt,
                     fifo_in_2_13_pt_V => fifo_in(2*NCALOFIFOS+13).pt,
                     fifo_in_2_14_pt_V => fifo_in(2*NCALOFIFOS+14).pt,
                     fifo_in_2_15_pt_V => fifo_in(2*NCALOFIFOS+15).pt,
                     fifo_in_2_16_pt_V => fifo_in(2*NCALOFIFOS+16).pt,
                     fifo_in_2_17_pt_V => fifo_in(2*NCALOFIFOS+17).pt,
                     fifo_in_2_18_pt_V => fifo_in(2*NCALOFIFOS+18).pt,
                     fifo_in_2_19_pt_V => fifo_in(2*NCALOFIFOS+19).pt,
                     fifo_in_0_0_eta_V  => fifo_in(0*NCALOFIFOS+ 0).eta,
                     fifo_in_0_1_eta_V  => fifo_in(0*NCALOFIFOS+ 1).eta,
                     fifo_in_0_2_eta_V  => fifo_in(0*NCALOFIFOS+ 2).eta,
                     fifo_in_0_3_eta_V  => fifo_in(0*NCALOFIFOS+ 3).eta,
                     fifo_in_0_4_eta_V  => fifo_in(0*NCALOFIFOS+ 4).eta,
                     fifo_in_0_5_eta_V  => fifo_in(0*NCALOFIFOS+ 5).eta,
                     fifo_in_0_6_eta_V  => fifo_in(0*NCALOFIFOS+ 6).eta,
                     fifo_in_0_7_eta_V  => fifo_in(0*NCALOFIFOS+ 7).eta,
                     fifo_in_0_8_eta_V  => fifo_in(0*NCALOFIFOS+ 8).eta,
                     fifo_in_0_9_eta_V  => fifo_in(0*NCALOFIFOS+ 9).eta,
                     fifo_in_0_10_eta_V => fifo_in(0*NCALOFIFOS+10).eta,
                     fifo_in_0_11_eta_V => fifo_in(0*NCALOFIFOS+11).eta,
                     fifo_in_0_12_eta_V => fifo_in(0*NCALOFIFOS+12).eta,
                     fifo_in_0_13_eta_V => fifo_in(0*NCALOFIFOS+13).eta,
                     fifo_in_0_14_eta_V => fifo_in(0*NCALOFIFOS+14).eta,
                     fifo_in_0_15_eta_V => fifo_in(0*NCALOFIFOS+15).eta,
                     fifo_in_0_16_eta_V => fifo_in(0*NCALOFIFOS+16).eta,
                     fifo_in_0_17_eta_V => fifo_in(0*NCALOFIFOS+17).eta,
                     fifo_in_0_18_eta_V => fifo_in(0*NCALOFIFOS+18).eta,
                     fifo_in_0_19_eta_V => fifo_in(0*NCALOFIFOS+19).eta,
                     fifo_in_1_0_eta_V  => fifo_in(1*NCALOFIFOS+ 0).eta,
                     fifo_in_1_1_eta_V  => fifo_in(1*NCALOFIFOS+ 1).eta,
                     fifo_in_1_2_eta_V  => fifo_in(1*NCALOFIFOS+ 2).eta,
                     fifo_in_1_3_eta_V  => fifo_in(1*NCALOFIFOS+ 3).eta,
                     fifo_in_1_4_eta_V  => fifo_in(1*NCALOFIFOS+ 4).eta,
                     fifo_in_1_5_eta_V  => fifo_in(1*NCALOFIFOS+ 5).eta,
                     fifo_in_1_6_eta_V  => fifo_in(1*NCALOFIFOS+ 6).eta,
                     fifo_in_1_7_eta_V  => fifo_in(1*NCALOFIFOS+ 7).eta,
                     fifo_in_1_8_eta_V  => fifo_in(1*NCALOFIFOS+ 8).eta,
                     fifo_in_1_9_eta_V  => fifo_in(1*NCALOFIFOS+ 9).eta,
                     fifo_in_1_10_eta_V => fifo_in(1*NCALOFIFOS+10).eta,
                     fifo_in_1_11_eta_V => fifo_in(1*NCALOFIFOS+11).eta,
                     fifo_in_1_12_eta_V => fifo_in(1*NCALOFIFOS+12).eta,
                     fifo_in_1_13_eta_V => fifo_in(1*NCALOFIFOS+13).eta,
                     fifo_in_1_14_eta_V => fifo_in(1*NCALOFIFOS+14).eta,
                     fifo_in_1_15_eta_V => fifo_in(1*NCALOFIFOS+15).eta,
                     fifo_in_1_16_eta_V => fifo_in(1*NCALOFIFOS+16).eta,
                     fifo_in_1_17_eta_V => fifo_in(1*NCALOFIFOS+17).eta,
                     fifo_in_1_18_eta_V => fifo_in(1*NCALOFIFOS+18).eta,
                     fifo_in_1_19_eta_V => fifo_in(1*NCALOFIFOS+19).eta,
                     fifo_in_2_0_eta_V  => fifo_in(2*NCALOFIFOS+ 0).eta,
                     fifo_in_2_1_eta_V  => fifo_in(2*NCALOFIFOS+ 1).eta,
                     fifo_in_2_2_eta_V  => fifo_in(2*NCALOFIFOS+ 2).eta,
                     fifo_in_2_3_eta_V  => fifo_in(2*NCALOFIFOS+ 3).eta,
                     fifo_in_2_4_eta_V  => fifo_in(2*NCALOFIFOS+ 4).eta,
                     fifo_in_2_5_eta_V  => fifo_in(2*NCALOFIFOS+ 5).eta,
                     fifo_in_2_6_eta_V  => fifo_in(2*NCALOFIFOS+ 6).eta,
                     fifo_in_2_7_eta_V  => fifo_in(2*NCALOFIFOS+ 7).eta,
                     fifo_in_2_8_eta_V  => fifo_in(2*NCALOFIFOS+ 8).eta,
                     fifo_in_2_9_eta_V  => fifo_in(2*NCALOFIFOS+ 9).eta,
                     fifo_in_2_10_eta_V => fifo_in(2*NCALOFIFOS+10).eta,
                     fifo_in_2_11_eta_V => fifo_in(2*NCALOFIFOS+11).eta,
                     fifo_in_2_12_eta_V => fifo_in(2*NCALOFIFOS+12).eta,
                     fifo_in_2_13_eta_V => fifo_in(2*NCALOFIFOS+13).eta,
                     fifo_in_2_14_eta_V => fifo_in(2*NCALOFIFOS+14).eta,
                     fifo_in_2_15_eta_V => fifo_in(2*NCALOFIFOS+15).eta,
                     fifo_in_2_16_eta_V => fifo_in(2*NCALOFIFOS+16).eta,
                     fifo_in_2_17_eta_V => fifo_in(2*NCALOFIFOS+17).eta,
                     fifo_in_2_18_eta_V => fifo_in(2*NCALOFIFOS+18).eta,
                     fifo_in_2_19_eta_V => fifo_in(2*NCALOFIFOS+19).eta,
                     fifo_in_0_0_phi_V  => fifo_in(0*NCALOFIFOS+ 0).phi,
                     fifo_in_0_1_phi_V  => fifo_in(0*NCALOFIFOS+ 1).phi,
                     fifo_in_0_2_phi_V  => fifo_in(0*NCALOFIFOS+ 2).phi,
                     fifo_in_0_3_phi_V  => fifo_in(0*NCALOFIFOS+ 3).phi,
                     fifo_in_0_4_phi_V  => fifo_in(0*NCALOFIFOS+ 4).phi,
                     fifo_in_0_5_phi_V  => fifo_in(0*NCALOFIFOS+ 5).phi,
                     fifo_in_0_6_phi_V  => fifo_in(0*NCALOFIFOS+ 6).phi,
                     fifo_in_0_7_phi_V  => fifo_in(0*NCALOFIFOS+ 7).phi,
                     fifo_in_0_8_phi_V  => fifo_in(0*NCALOFIFOS+ 8).phi,
                     fifo_in_0_9_phi_V  => fifo_in(0*NCALOFIFOS+ 9).phi,
                     fifo_in_0_10_phi_V => fifo_in(0*NCALOFIFOS+10).phi,
                     fifo_in_0_11_phi_V => fifo_in(0*NCALOFIFOS+11).phi,
                     fifo_in_0_12_phi_V => fifo_in(0*NCALOFIFOS+12).phi,
                     fifo_in_0_13_phi_V => fifo_in(0*NCALOFIFOS+13).phi,
                     fifo_in_0_14_phi_V => fifo_in(0*NCALOFIFOS+14).phi,
                     fifo_in_0_15_phi_V => fifo_in(0*NCALOFIFOS+15).phi,
                     fifo_in_0_16_phi_V => fifo_in(0*NCALOFIFOS+16).phi,
                     fifo_in_0_17_phi_V => fifo_in(0*NCALOFIFOS+17).phi,
                     fifo_in_0_18_phi_V => fifo_in(0*NCALOFIFOS+18).phi,
                     fifo_in_0_19_phi_V => fifo_in(0*NCALOFIFOS+19).phi,
                     fifo_in_1_0_phi_V  => fifo_in(1*NCALOFIFOS+ 0).phi,
                     fifo_in_1_1_phi_V  => fifo_in(1*NCALOFIFOS+ 1).phi,
                     fifo_in_1_2_phi_V  => fifo_in(1*NCALOFIFOS+ 2).phi,
                     fifo_in_1_3_phi_V  => fifo_in(1*NCALOFIFOS+ 3).phi,
                     fifo_in_1_4_phi_V  => fifo_in(1*NCALOFIFOS+ 4).phi,
                     fifo_in_1_5_phi_V  => fifo_in(1*NCALOFIFOS+ 5).phi,
                     fifo_in_1_6_phi_V  => fifo_in(1*NCALOFIFOS+ 6).phi,
                     fifo_in_1_7_phi_V  => fifo_in(1*NCALOFIFOS+ 7).phi,
                     fifo_in_1_8_phi_V  => fifo_in(1*NCALOFIFOS+ 8).phi,
                     fifo_in_1_9_phi_V  => fifo_in(1*NCALOFIFOS+ 9).phi,
                     fifo_in_1_10_phi_V => fifo_in(1*NCALOFIFOS+10).phi,
                     fifo_in_1_11_phi_V => fifo_in(1*NCALOFIFOS+11).phi,
                     fifo_in_1_12_phi_V => fifo_in(1*NCALOFIFOS+12).phi,
                     fifo_in_1_13_phi_V => fifo_in(1*NCALOFIFOS+13).phi,
                     fifo_in_1_14_phi_V => fifo_in(1*NCALOFIFOS+14).phi,
                     fifo_in_1_15_phi_V => fifo_in(1*NCALOFIFOS+15).phi,
                     fifo_in_1_16_phi_V => fifo_in(1*NCALOFIFOS+16).phi,
                     fifo_in_1_17_phi_V => fifo_in(1*NCALOFIFOS+17).phi,
                     fifo_in_1_18_phi_V => fifo_in(1*NCALOFIFOS+18).phi,
                     fifo_in_1_19_phi_V => fifo_in(1*NCALOFIFOS+19).phi,
                     fifo_in_2_0_phi_V  => fifo_in(2*NCALOFIFOS+ 0).phi,
                     fifo_in_2_1_phi_V  => fifo_in(2*NCALOFIFOS+ 1).phi,
                     fifo_in_2_2_phi_V  => fifo_in(2*NCALOFIFOS+ 2).phi,
                     fifo_in_2_3_phi_V  => fifo_in(2*NCALOFIFOS+ 3).phi,
                     fifo_in_2_4_phi_V  => fifo_in(2*NCALOFIFOS+ 4).phi,
                     fifo_in_2_5_phi_V  => fifo_in(2*NCALOFIFOS+ 5).phi,
                     fifo_in_2_6_phi_V  => fifo_in(2*NCALOFIFOS+ 6).phi,
                     fifo_in_2_7_phi_V  => fifo_in(2*NCALOFIFOS+ 7).phi,
                     fifo_in_2_8_phi_V  => fifo_in(2*NCALOFIFOS+ 8).phi,
                     fifo_in_2_9_phi_V  => fifo_in(2*NCALOFIFOS+ 9).phi,
                     fifo_in_2_10_phi_V => fifo_in(2*NCALOFIFOS+10).phi,
                     fifo_in_2_11_phi_V => fifo_in(2*NCALOFIFOS+11).phi,
                     fifo_in_2_12_phi_V => fifo_in(2*NCALOFIFOS+12).phi,
                     fifo_in_2_13_phi_V => fifo_in(2*NCALOFIFOS+13).phi,
                     fifo_in_2_14_phi_V => fifo_in(2*NCALOFIFOS+14).phi,
                     fifo_in_2_15_phi_V => fifo_in(2*NCALOFIFOS+15).phi,
                     fifo_in_2_16_phi_V => fifo_in(2*NCALOFIFOS+16).phi,
                     fifo_in_2_17_phi_V => fifo_in(2*NCALOFIFOS+17).phi,
                     fifo_in_2_18_phi_V => fifo_in(2*NCALOFIFOS+18).phi,
                     fifo_in_2_19_phi_V => fifo_in(2*NCALOFIFOS+19).phi,
                     fifo_in_0_0_rest_V  => fifo_in(0*NCALOFIFOS+ 0).rest,
                     fifo_in_0_1_rest_V  => fifo_in(0*NCALOFIFOS+ 1).rest,
                     fifo_in_0_2_rest_V  => fifo_in(0*NCALOFIFOS+ 2).rest,
                     fifo_in_0_3_rest_V  => fifo_in(0*NCALOFIFOS+ 3).rest,
                     fifo_in_0_4_rest_V  => fifo_in(0*NCALOFIFOS+ 4).rest,
                     fifo_in_0_5_rest_V  => fifo_in(0*NCALOFIFOS+ 5).rest,
                     fifo_in_0_6_rest_V  => fifo_in(0*NCALOFIFOS+ 6).rest,
                     fifo_in_0_7_rest_V  => fifo_in(0*NCALOFIFOS+ 7).rest,
                     fifo_in_0_8_rest_V  => fifo_in(0*NCALOFIFOS+ 8).rest,
                     fifo_in_0_9_rest_V  => fifo_in(0*NCALOFIFOS+ 9).rest,
                     fifo_in_0_10_rest_V => fifo_in(0*NCALOFIFOS+10).rest,
                     fifo_in_0_11_rest_V => fifo_in(0*NCALOFIFOS+11).rest,
                     fifo_in_0_12_rest_V => fifo_in(0*NCALOFIFOS+12).rest,
                     fifo_in_0_13_rest_V => fifo_in(0*NCALOFIFOS+13).rest,
                     fifo_in_0_14_rest_V => fifo_in(0*NCALOFIFOS+14).rest,
                     fifo_in_0_15_rest_V => fifo_in(0*NCALOFIFOS+15).rest,
                     fifo_in_0_16_rest_V => fifo_in(0*NCALOFIFOS+16).rest,
                     fifo_in_0_17_rest_V => fifo_in(0*NCALOFIFOS+17).rest,
                     fifo_in_0_18_rest_V => fifo_in(0*NCALOFIFOS+18).rest,
                     fifo_in_0_19_rest_V => fifo_in(0*NCALOFIFOS+19).rest,
                     fifo_in_1_0_rest_V  => fifo_in(1*NCALOFIFOS+ 0).rest,
                     fifo_in_1_1_rest_V  => fifo_in(1*NCALOFIFOS+ 1).rest,
                     fifo_in_1_2_rest_V  => fifo_in(1*NCALOFIFOS+ 2).rest,
                     fifo_in_1_3_rest_V  => fifo_in(1*NCALOFIFOS+ 3).rest,
                     fifo_in_1_4_rest_V  => fifo_in(1*NCALOFIFOS+ 4).rest,
                     fifo_in_1_5_rest_V  => fifo_in(1*NCALOFIFOS+ 5).rest,
                     fifo_in_1_6_rest_V  => fifo_in(1*NCALOFIFOS+ 6).rest,
                     fifo_in_1_7_rest_V  => fifo_in(1*NCALOFIFOS+ 7).rest,
                     fifo_in_1_8_rest_V  => fifo_in(1*NCALOFIFOS+ 8).rest,
                     fifo_in_1_9_rest_V  => fifo_in(1*NCALOFIFOS+ 9).rest,
                     fifo_in_1_10_rest_V => fifo_in(1*NCALOFIFOS+10).rest,
                     fifo_in_1_11_rest_V => fifo_in(1*NCALOFIFOS+11).rest,
                     fifo_in_1_12_rest_V => fifo_in(1*NCALOFIFOS+12).rest,
                     fifo_in_1_13_rest_V => fifo_in(1*NCALOFIFOS+13).rest,
                     fifo_in_1_14_rest_V => fifo_in(1*NCALOFIFOS+14).rest,
                     fifo_in_1_15_rest_V => fifo_in(1*NCALOFIFOS+15).rest,
                     fifo_in_1_16_rest_V => fifo_in(1*NCALOFIFOS+16).rest,
                     fifo_in_1_17_rest_V => fifo_in(1*NCALOFIFOS+17).rest,
                     fifo_in_1_18_rest_V => fifo_in(1*NCALOFIFOS+18).rest,
                     fifo_in_1_19_rest_V => fifo_in(1*NCALOFIFOS+19).rest,
                     fifo_in_2_0_rest_V  => fifo_in(2*NCALOFIFOS+ 0).rest,
                     fifo_in_2_1_rest_V  => fifo_in(2*NCALOFIFOS+ 1).rest,
                     fifo_in_2_2_rest_V  => fifo_in(2*NCALOFIFOS+ 2).rest,
                     fifo_in_2_3_rest_V  => fifo_in(2*NCALOFIFOS+ 3).rest,
                     fifo_in_2_4_rest_V  => fifo_in(2*NCALOFIFOS+ 4).rest,
                     fifo_in_2_5_rest_V  => fifo_in(2*NCALOFIFOS+ 5).rest,
                     fifo_in_2_6_rest_V  => fifo_in(2*NCALOFIFOS+ 6).rest,
                     fifo_in_2_7_rest_V  => fifo_in(2*NCALOFIFOS+ 7).rest,
                     fifo_in_2_8_rest_V  => fifo_in(2*NCALOFIFOS+ 8).rest,
                     fifo_in_2_9_rest_V  => fifo_in(2*NCALOFIFOS+ 9).rest,
                     fifo_in_2_10_rest_V => fifo_in(2*NCALOFIFOS+10).rest,
                     fifo_in_2_11_rest_V => fifo_in(2*NCALOFIFOS+11).rest,
                     fifo_in_2_12_rest_V => fifo_in(2*NCALOFIFOS+12).rest,
                     fifo_in_2_13_rest_V => fifo_in(2*NCALOFIFOS+13).rest,
                     fifo_in_2_14_rest_V => fifo_in(2*NCALOFIFOS+14).rest,
                     fifo_in_2_15_rest_V => fifo_in(2*NCALOFIFOS+15).rest,
                     fifo_in_2_16_rest_V => fifo_in(2*NCALOFIFOS+16).rest,
                     fifo_in_2_17_rest_V => fifo_in(2*NCALOFIFOS+17).rest,
                     fifo_in_2_18_rest_V => fifo_in(2*NCALOFIFOS+18).rest,
                     fifo_in_2_19_rest_V => fifo_in(2*NCALOFIFOS+19).rest,
                     fifo_write_0_0  => fifo_write(0*NCALOFIFOS+ 0),
                     fifo_write_0_1  => fifo_write(0*NCALOFIFOS+ 1),
                     fifo_write_0_2  => fifo_write(0*NCALOFIFOS+ 2),
                     fifo_write_0_3  => fifo_write(0*NCALOFIFOS+ 3),
                     fifo_write_0_4  => fifo_write(0*NCALOFIFOS+ 4),
                     fifo_write_0_5  => fifo_write(0*NCALOFIFOS+ 5),
                     fifo_write_0_6  => fifo_write(0*NCALOFIFOS+ 6),
                     fifo_write_0_7  => fifo_write(0*NCALOFIFOS+ 7),
                     fifo_write_0_8  => fifo_write(0*NCALOFIFOS+ 8),
                     fifo_write_0_9  => fifo_write(0*NCALOFIFOS+ 9),
                     fifo_write_0_10 => fifo_write(0*NCALOFIFOS+10),
                     fifo_write_0_11 => fifo_write(0*NCALOFIFOS+11),
                     fifo_write_0_12 => fifo_write(0*NCALOFIFOS+12),
                     fifo_write_0_13 => fifo_write(0*NCALOFIFOS+13),
                     fifo_write_0_14 => fifo_write(0*NCALOFIFOS+14),
                     fifo_write_0_15 => fifo_write(0*NCALOFIFOS+15),
                     fifo_write_0_16 => fifo_write(0*NCALOFIFOS+16),
                     fifo_write_0_17 => fifo_write(0*NCALOFIFOS+17),
                     fifo_write_0_18 => fifo_write(0*NCALOFIFOS+18),
                     fifo_write_0_19 => fifo_write(0*NCALOFIFOS+19),
                     fifo_write_1_0  => fifo_write(1*NCALOFIFOS+ 0),
                     fifo_write_1_1  => fifo_write(1*NCALOFIFOS+ 1),
                     fifo_write_1_2  => fifo_write(1*NCALOFIFOS+ 2),
                     fifo_write_1_3  => fifo_write(1*NCALOFIFOS+ 3),
                     fifo_write_1_4  => fifo_write(1*NCALOFIFOS+ 4),
                     fifo_write_1_5  => fifo_write(1*NCALOFIFOS+ 5),
                     fifo_write_1_6  => fifo_write(1*NCALOFIFOS+ 6),
                     fifo_write_1_7  => fifo_write(1*NCALOFIFOS+ 7),
                     fifo_write_1_8  => fifo_write(1*NCALOFIFOS+ 8),
                     fifo_write_1_9  => fifo_write(1*NCALOFIFOS+ 9),
                     fifo_write_1_10 => fifo_write(1*NCALOFIFOS+10),
                     fifo_write_1_11 => fifo_write(1*NCALOFIFOS+11),
                     fifo_write_1_12 => fifo_write(1*NCALOFIFOS+12),
                     fifo_write_1_13 => fifo_write(1*NCALOFIFOS+13),
                     fifo_write_1_14 => fifo_write(1*NCALOFIFOS+14),
                     fifo_write_1_15 => fifo_write(1*NCALOFIFOS+15),
                     fifo_write_1_16 => fifo_write(1*NCALOFIFOS+16),
                     fifo_write_1_17 => fifo_write(1*NCALOFIFOS+17),
                     fifo_write_1_18 => fifo_write(1*NCALOFIFOS+18),
                     fifo_write_1_19 => fifo_write(1*NCALOFIFOS+19),
                     fifo_write_2_0  => fifo_write(2*NCALOFIFOS+ 0),
                     fifo_write_2_1  => fifo_write(2*NCALOFIFOS+ 1),
                     fifo_write_2_2  => fifo_write(2*NCALOFIFOS+ 2),
                     fifo_write_2_3  => fifo_write(2*NCALOFIFOS+ 3),
                     fifo_write_2_4  => fifo_write(2*NCALOFIFOS+ 4),
                     fifo_write_2_5  => fifo_write(2*NCALOFIFOS+ 5),
                     fifo_write_2_6  => fifo_write(2*NCALOFIFOS+ 6),
                     fifo_write_2_7  => fifo_write(2*NCALOFIFOS+ 7),
                     fifo_write_2_8  => fifo_write(2*NCALOFIFOS+ 8),
                     fifo_write_2_9  => fifo_write(2*NCALOFIFOS+ 9),
                     fifo_write_2_10 => fifo_write(2*NCALOFIFOS+10),
                     fifo_write_2_11 => fifo_write(2*NCALOFIFOS+11),
                     fifo_write_2_12 => fifo_write(2*NCALOFIFOS+12),
                     fifo_write_2_13 => fifo_write(2*NCALOFIFOS+13),
                     fifo_write_2_14 => fifo_write(2*NCALOFIFOS+14),
                     fifo_write_2_15 => fifo_write(2*NCALOFIFOS+15),
                     fifo_write_2_16 => fifo_write(2*NCALOFIFOS+16),
                     fifo_write_2_17 => fifo_write(2*NCALOFIFOS+17),
                     fifo_write_2_18 => fifo_write(2*NCALOFIFOS+18),
                     fifo_write_2_19 => fifo_write(2*NCALOFIFOS+19)
                 );

    fifo_slice : entity work.calo_router_fifo_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     newevent => newevent_del,
                     fifo_in_0_0_pt_V  => fifo_in(0*NCALOFIFOS+ 0).pt,
                     fifo_in_0_1_pt_V  => fifo_in(0*NCALOFIFOS+ 1).pt,
                     fifo_in_0_2_pt_V  => fifo_in(0*NCALOFIFOS+ 2).pt,
                     fifo_in_0_3_pt_V  => fifo_in(0*NCALOFIFOS+ 3).pt,
                     fifo_in_0_4_pt_V  => fifo_in(0*NCALOFIFOS+ 4).pt,
                     fifo_in_0_5_pt_V  => fifo_in(0*NCALOFIFOS+ 5).pt,
                     fifo_in_0_6_pt_V  => fifo_in(0*NCALOFIFOS+ 6).pt,
                     fifo_in_0_7_pt_V  => fifo_in(0*NCALOFIFOS+ 7).pt,
                     fifo_in_0_8_pt_V  => fifo_in(0*NCALOFIFOS+ 8).pt,
                     fifo_in_0_9_pt_V  => fifo_in(0*NCALOFIFOS+ 9).pt,
                     fifo_in_0_10_pt_V => fifo_in(0*NCALOFIFOS+10).pt,
                     fifo_in_0_11_pt_V => fifo_in(0*NCALOFIFOS+11).pt,
                     fifo_in_0_12_pt_V => fifo_in(0*NCALOFIFOS+12).pt,
                     fifo_in_0_13_pt_V => fifo_in(0*NCALOFIFOS+13).pt,
                     fifo_in_0_14_pt_V => fifo_in(0*NCALOFIFOS+14).pt,
                     fifo_in_0_15_pt_V => fifo_in(0*NCALOFIFOS+15).pt,
                     fifo_in_0_16_pt_V => fifo_in(0*NCALOFIFOS+16).pt,
                     fifo_in_0_17_pt_V => fifo_in(0*NCALOFIFOS+17).pt,
                     fifo_in_0_18_pt_V => fifo_in(0*NCALOFIFOS+18).pt,
                     fifo_in_0_19_pt_V => fifo_in(0*NCALOFIFOS+19).pt,
                     fifo_in_1_0_pt_V  => fifo_in(1*NCALOFIFOS+ 0).pt,
                     fifo_in_1_1_pt_V  => fifo_in(1*NCALOFIFOS+ 1).pt,
                     fifo_in_1_2_pt_V  => fifo_in(1*NCALOFIFOS+ 2).pt,
                     fifo_in_1_3_pt_V  => fifo_in(1*NCALOFIFOS+ 3).pt,
                     fifo_in_1_4_pt_V  => fifo_in(1*NCALOFIFOS+ 4).pt,
                     fifo_in_1_5_pt_V  => fifo_in(1*NCALOFIFOS+ 5).pt,
                     fifo_in_1_6_pt_V  => fifo_in(1*NCALOFIFOS+ 6).pt,
                     fifo_in_1_7_pt_V  => fifo_in(1*NCALOFIFOS+ 7).pt,
                     fifo_in_1_8_pt_V  => fifo_in(1*NCALOFIFOS+ 8).pt,
                     fifo_in_1_9_pt_V  => fifo_in(1*NCALOFIFOS+ 9).pt,
                     fifo_in_1_10_pt_V => fifo_in(1*NCALOFIFOS+10).pt,
                     fifo_in_1_11_pt_V => fifo_in(1*NCALOFIFOS+11).pt,
                     fifo_in_1_12_pt_V => fifo_in(1*NCALOFIFOS+12).pt,
                     fifo_in_1_13_pt_V => fifo_in(1*NCALOFIFOS+13).pt,
                     fifo_in_1_14_pt_V => fifo_in(1*NCALOFIFOS+14).pt,
                     fifo_in_1_15_pt_V => fifo_in(1*NCALOFIFOS+15).pt,
                     fifo_in_1_16_pt_V => fifo_in(1*NCALOFIFOS+16).pt,
                     fifo_in_1_17_pt_V => fifo_in(1*NCALOFIFOS+17).pt,
                     fifo_in_1_18_pt_V => fifo_in(1*NCALOFIFOS+18).pt,
                     fifo_in_1_19_pt_V => fifo_in(1*NCALOFIFOS+19).pt,
                     fifo_in_2_0_pt_V  => fifo_in(2*NCALOFIFOS+ 0).pt,
                     fifo_in_2_1_pt_V  => fifo_in(2*NCALOFIFOS+ 1).pt,
                     fifo_in_2_2_pt_V  => fifo_in(2*NCALOFIFOS+ 2).pt,
                     fifo_in_2_3_pt_V  => fifo_in(2*NCALOFIFOS+ 3).pt,
                     fifo_in_2_4_pt_V  => fifo_in(2*NCALOFIFOS+ 4).pt,
                     fifo_in_2_5_pt_V  => fifo_in(2*NCALOFIFOS+ 5).pt,
                     fifo_in_2_6_pt_V  => fifo_in(2*NCALOFIFOS+ 6).pt,
                     fifo_in_2_7_pt_V  => fifo_in(2*NCALOFIFOS+ 7).pt,
                     fifo_in_2_8_pt_V  => fifo_in(2*NCALOFIFOS+ 8).pt,
                     fifo_in_2_9_pt_V  => fifo_in(2*NCALOFIFOS+ 9).pt,
                     fifo_in_2_10_pt_V => fifo_in(2*NCALOFIFOS+10).pt,
                     fifo_in_2_11_pt_V => fifo_in(2*NCALOFIFOS+11).pt,
                     fifo_in_2_12_pt_V => fifo_in(2*NCALOFIFOS+12).pt,
                     fifo_in_2_13_pt_V => fifo_in(2*NCALOFIFOS+13).pt,
                     fifo_in_2_14_pt_V => fifo_in(2*NCALOFIFOS+14).pt,
                     fifo_in_2_15_pt_V => fifo_in(2*NCALOFIFOS+15).pt,
                     fifo_in_2_16_pt_V => fifo_in(2*NCALOFIFOS+16).pt,
                     fifo_in_2_17_pt_V => fifo_in(2*NCALOFIFOS+17).pt,
                     fifo_in_2_18_pt_V => fifo_in(2*NCALOFIFOS+18).pt,
                     fifo_in_2_19_pt_V => fifo_in(2*NCALOFIFOS+19).pt,
                     fifo_in_0_0_eta_V  => fifo_in(0*NCALOFIFOS+ 0).eta,
                     fifo_in_0_1_eta_V  => fifo_in(0*NCALOFIFOS+ 1).eta,
                     fifo_in_0_2_eta_V  => fifo_in(0*NCALOFIFOS+ 2).eta,
                     fifo_in_0_3_eta_V  => fifo_in(0*NCALOFIFOS+ 3).eta,
                     fifo_in_0_4_eta_V  => fifo_in(0*NCALOFIFOS+ 4).eta,
                     fifo_in_0_5_eta_V  => fifo_in(0*NCALOFIFOS+ 5).eta,
                     fifo_in_0_6_eta_V  => fifo_in(0*NCALOFIFOS+ 6).eta,
                     fifo_in_0_7_eta_V  => fifo_in(0*NCALOFIFOS+ 7).eta,
                     fifo_in_0_8_eta_V  => fifo_in(0*NCALOFIFOS+ 8).eta,
                     fifo_in_0_9_eta_V  => fifo_in(0*NCALOFIFOS+ 9).eta,
                     fifo_in_0_10_eta_V => fifo_in(0*NCALOFIFOS+10).eta,
                     fifo_in_0_11_eta_V => fifo_in(0*NCALOFIFOS+11).eta,
                     fifo_in_0_12_eta_V => fifo_in(0*NCALOFIFOS+12).eta,
                     fifo_in_0_13_eta_V => fifo_in(0*NCALOFIFOS+13).eta,
                     fifo_in_0_14_eta_V => fifo_in(0*NCALOFIFOS+14).eta,
                     fifo_in_0_15_eta_V => fifo_in(0*NCALOFIFOS+15).eta,
                     fifo_in_0_16_eta_V => fifo_in(0*NCALOFIFOS+16).eta,
                     fifo_in_0_17_eta_V => fifo_in(0*NCALOFIFOS+17).eta,
                     fifo_in_0_18_eta_V => fifo_in(0*NCALOFIFOS+18).eta,
                     fifo_in_0_19_eta_V => fifo_in(0*NCALOFIFOS+19).eta,
                     fifo_in_1_0_eta_V  => fifo_in(1*NCALOFIFOS+ 0).eta,
                     fifo_in_1_1_eta_V  => fifo_in(1*NCALOFIFOS+ 1).eta,
                     fifo_in_1_2_eta_V  => fifo_in(1*NCALOFIFOS+ 2).eta,
                     fifo_in_1_3_eta_V  => fifo_in(1*NCALOFIFOS+ 3).eta,
                     fifo_in_1_4_eta_V  => fifo_in(1*NCALOFIFOS+ 4).eta,
                     fifo_in_1_5_eta_V  => fifo_in(1*NCALOFIFOS+ 5).eta,
                     fifo_in_1_6_eta_V  => fifo_in(1*NCALOFIFOS+ 6).eta,
                     fifo_in_1_7_eta_V  => fifo_in(1*NCALOFIFOS+ 7).eta,
                     fifo_in_1_8_eta_V  => fifo_in(1*NCALOFIFOS+ 8).eta,
                     fifo_in_1_9_eta_V  => fifo_in(1*NCALOFIFOS+ 9).eta,
                     fifo_in_1_10_eta_V => fifo_in(1*NCALOFIFOS+10).eta,
                     fifo_in_1_11_eta_V => fifo_in(1*NCALOFIFOS+11).eta,
                     fifo_in_1_12_eta_V => fifo_in(1*NCALOFIFOS+12).eta,
                     fifo_in_1_13_eta_V => fifo_in(1*NCALOFIFOS+13).eta,
                     fifo_in_1_14_eta_V => fifo_in(1*NCALOFIFOS+14).eta,
                     fifo_in_1_15_eta_V => fifo_in(1*NCALOFIFOS+15).eta,
                     fifo_in_1_16_eta_V => fifo_in(1*NCALOFIFOS+16).eta,
                     fifo_in_1_17_eta_V => fifo_in(1*NCALOFIFOS+17).eta,
                     fifo_in_1_18_eta_V => fifo_in(1*NCALOFIFOS+18).eta,
                     fifo_in_1_19_eta_V => fifo_in(1*NCALOFIFOS+19).eta,
                     fifo_in_2_0_eta_V  => fifo_in(2*NCALOFIFOS+ 0).eta,
                     fifo_in_2_1_eta_V  => fifo_in(2*NCALOFIFOS+ 1).eta,
                     fifo_in_2_2_eta_V  => fifo_in(2*NCALOFIFOS+ 2).eta,
                     fifo_in_2_3_eta_V  => fifo_in(2*NCALOFIFOS+ 3).eta,
                     fifo_in_2_4_eta_V  => fifo_in(2*NCALOFIFOS+ 4).eta,
                     fifo_in_2_5_eta_V  => fifo_in(2*NCALOFIFOS+ 5).eta,
                     fifo_in_2_6_eta_V  => fifo_in(2*NCALOFIFOS+ 6).eta,
                     fifo_in_2_7_eta_V  => fifo_in(2*NCALOFIFOS+ 7).eta,
                     fifo_in_2_8_eta_V  => fifo_in(2*NCALOFIFOS+ 8).eta,
                     fifo_in_2_9_eta_V  => fifo_in(2*NCALOFIFOS+ 9).eta,
                     fifo_in_2_10_eta_V => fifo_in(2*NCALOFIFOS+10).eta,
                     fifo_in_2_11_eta_V => fifo_in(2*NCALOFIFOS+11).eta,
                     fifo_in_2_12_eta_V => fifo_in(2*NCALOFIFOS+12).eta,
                     fifo_in_2_13_eta_V => fifo_in(2*NCALOFIFOS+13).eta,
                     fifo_in_2_14_eta_V => fifo_in(2*NCALOFIFOS+14).eta,
                     fifo_in_2_15_eta_V => fifo_in(2*NCALOFIFOS+15).eta,
                     fifo_in_2_16_eta_V => fifo_in(2*NCALOFIFOS+16).eta,
                     fifo_in_2_17_eta_V => fifo_in(2*NCALOFIFOS+17).eta,
                     fifo_in_2_18_eta_V => fifo_in(2*NCALOFIFOS+18).eta,
                     fifo_in_2_19_eta_V => fifo_in(2*NCALOFIFOS+19).eta,
                     fifo_in_0_0_phi_V  => fifo_in(0*NCALOFIFOS+ 0).phi,
                     fifo_in_0_1_phi_V  => fifo_in(0*NCALOFIFOS+ 1).phi,
                     fifo_in_0_2_phi_V  => fifo_in(0*NCALOFIFOS+ 2).phi,
                     fifo_in_0_3_phi_V  => fifo_in(0*NCALOFIFOS+ 3).phi,
                     fifo_in_0_4_phi_V  => fifo_in(0*NCALOFIFOS+ 4).phi,
                     fifo_in_0_5_phi_V  => fifo_in(0*NCALOFIFOS+ 5).phi,
                     fifo_in_0_6_phi_V  => fifo_in(0*NCALOFIFOS+ 6).phi,
                     fifo_in_0_7_phi_V  => fifo_in(0*NCALOFIFOS+ 7).phi,
                     fifo_in_0_8_phi_V  => fifo_in(0*NCALOFIFOS+ 8).phi,
                     fifo_in_0_9_phi_V  => fifo_in(0*NCALOFIFOS+ 9).phi,
                     fifo_in_0_10_phi_V => fifo_in(0*NCALOFIFOS+10).phi,
                     fifo_in_0_11_phi_V => fifo_in(0*NCALOFIFOS+11).phi,
                     fifo_in_0_12_phi_V => fifo_in(0*NCALOFIFOS+12).phi,
                     fifo_in_0_13_phi_V => fifo_in(0*NCALOFIFOS+13).phi,
                     fifo_in_0_14_phi_V => fifo_in(0*NCALOFIFOS+14).phi,
                     fifo_in_0_15_phi_V => fifo_in(0*NCALOFIFOS+15).phi,
                     fifo_in_0_16_phi_V => fifo_in(0*NCALOFIFOS+16).phi,
                     fifo_in_0_17_phi_V => fifo_in(0*NCALOFIFOS+17).phi,
                     fifo_in_0_18_phi_V => fifo_in(0*NCALOFIFOS+18).phi,
                     fifo_in_0_19_phi_V => fifo_in(0*NCALOFIFOS+19).phi,
                     fifo_in_1_0_phi_V  => fifo_in(1*NCALOFIFOS+ 0).phi,
                     fifo_in_1_1_phi_V  => fifo_in(1*NCALOFIFOS+ 1).phi,
                     fifo_in_1_2_phi_V  => fifo_in(1*NCALOFIFOS+ 2).phi,
                     fifo_in_1_3_phi_V  => fifo_in(1*NCALOFIFOS+ 3).phi,
                     fifo_in_1_4_phi_V  => fifo_in(1*NCALOFIFOS+ 4).phi,
                     fifo_in_1_5_phi_V  => fifo_in(1*NCALOFIFOS+ 5).phi,
                     fifo_in_1_6_phi_V  => fifo_in(1*NCALOFIFOS+ 6).phi,
                     fifo_in_1_7_phi_V  => fifo_in(1*NCALOFIFOS+ 7).phi,
                     fifo_in_1_8_phi_V  => fifo_in(1*NCALOFIFOS+ 8).phi,
                     fifo_in_1_9_phi_V  => fifo_in(1*NCALOFIFOS+ 9).phi,
                     fifo_in_1_10_phi_V => fifo_in(1*NCALOFIFOS+10).phi,
                     fifo_in_1_11_phi_V => fifo_in(1*NCALOFIFOS+11).phi,
                     fifo_in_1_12_phi_V => fifo_in(1*NCALOFIFOS+12).phi,
                     fifo_in_1_13_phi_V => fifo_in(1*NCALOFIFOS+13).phi,
                     fifo_in_1_14_phi_V => fifo_in(1*NCALOFIFOS+14).phi,
                     fifo_in_1_15_phi_V => fifo_in(1*NCALOFIFOS+15).phi,
                     fifo_in_1_16_phi_V => fifo_in(1*NCALOFIFOS+16).phi,
                     fifo_in_1_17_phi_V => fifo_in(1*NCALOFIFOS+17).phi,
                     fifo_in_1_18_phi_V => fifo_in(1*NCALOFIFOS+18).phi,
                     fifo_in_1_19_phi_V => fifo_in(1*NCALOFIFOS+19).phi,
                     fifo_in_2_0_phi_V  => fifo_in(2*NCALOFIFOS+ 0).phi,
                     fifo_in_2_1_phi_V  => fifo_in(2*NCALOFIFOS+ 1).phi,
                     fifo_in_2_2_phi_V  => fifo_in(2*NCALOFIFOS+ 2).phi,
                     fifo_in_2_3_phi_V  => fifo_in(2*NCALOFIFOS+ 3).phi,
                     fifo_in_2_4_phi_V  => fifo_in(2*NCALOFIFOS+ 4).phi,
                     fifo_in_2_5_phi_V  => fifo_in(2*NCALOFIFOS+ 5).phi,
                     fifo_in_2_6_phi_V  => fifo_in(2*NCALOFIFOS+ 6).phi,
                     fifo_in_2_7_phi_V  => fifo_in(2*NCALOFIFOS+ 7).phi,
                     fifo_in_2_8_phi_V  => fifo_in(2*NCALOFIFOS+ 8).phi,
                     fifo_in_2_9_phi_V  => fifo_in(2*NCALOFIFOS+ 9).phi,
                     fifo_in_2_10_phi_V => fifo_in(2*NCALOFIFOS+10).phi,
                     fifo_in_2_11_phi_V => fifo_in(2*NCALOFIFOS+11).phi,
                     fifo_in_2_12_phi_V => fifo_in(2*NCALOFIFOS+12).phi,
                     fifo_in_2_13_phi_V => fifo_in(2*NCALOFIFOS+13).phi,
                     fifo_in_2_14_phi_V => fifo_in(2*NCALOFIFOS+14).phi,
                     fifo_in_2_15_phi_V => fifo_in(2*NCALOFIFOS+15).phi,
                     fifo_in_2_16_phi_V => fifo_in(2*NCALOFIFOS+16).phi,
                     fifo_in_2_17_phi_V => fifo_in(2*NCALOFIFOS+17).phi,
                     fifo_in_2_18_phi_V => fifo_in(2*NCALOFIFOS+18).phi,
                     fifo_in_2_19_phi_V => fifo_in(2*NCALOFIFOS+19).phi,
                     fifo_in_0_0_rest_V  => fifo_in(0*NCALOFIFOS+ 0).rest,
                     fifo_in_0_1_rest_V  => fifo_in(0*NCALOFIFOS+ 1).rest,
                     fifo_in_0_2_rest_V  => fifo_in(0*NCALOFIFOS+ 2).rest,
                     fifo_in_0_3_rest_V  => fifo_in(0*NCALOFIFOS+ 3).rest,
                     fifo_in_0_4_rest_V  => fifo_in(0*NCALOFIFOS+ 4).rest,
                     fifo_in_0_5_rest_V  => fifo_in(0*NCALOFIFOS+ 5).rest,
                     fifo_in_0_6_rest_V  => fifo_in(0*NCALOFIFOS+ 6).rest,
                     fifo_in_0_7_rest_V  => fifo_in(0*NCALOFIFOS+ 7).rest,
                     fifo_in_0_8_rest_V  => fifo_in(0*NCALOFIFOS+ 8).rest,
                     fifo_in_0_9_rest_V  => fifo_in(0*NCALOFIFOS+ 9).rest,
                     fifo_in_0_10_rest_V => fifo_in(0*NCALOFIFOS+10).rest,
                     fifo_in_0_11_rest_V => fifo_in(0*NCALOFIFOS+11).rest,
                     fifo_in_0_12_rest_V => fifo_in(0*NCALOFIFOS+12).rest,
                     fifo_in_0_13_rest_V => fifo_in(0*NCALOFIFOS+13).rest,
                     fifo_in_0_14_rest_V => fifo_in(0*NCALOFIFOS+14).rest,
                     fifo_in_0_15_rest_V => fifo_in(0*NCALOFIFOS+15).rest,
                     fifo_in_0_16_rest_V => fifo_in(0*NCALOFIFOS+16).rest,
                     fifo_in_0_17_rest_V => fifo_in(0*NCALOFIFOS+17).rest,
                     fifo_in_0_18_rest_V => fifo_in(0*NCALOFIFOS+18).rest,
                     fifo_in_0_19_rest_V => fifo_in(0*NCALOFIFOS+19).rest,
                     fifo_in_1_0_rest_V  => fifo_in(1*NCALOFIFOS+ 0).rest,
                     fifo_in_1_1_rest_V  => fifo_in(1*NCALOFIFOS+ 1).rest,
                     fifo_in_1_2_rest_V  => fifo_in(1*NCALOFIFOS+ 2).rest,
                     fifo_in_1_3_rest_V  => fifo_in(1*NCALOFIFOS+ 3).rest,
                     fifo_in_1_4_rest_V  => fifo_in(1*NCALOFIFOS+ 4).rest,
                     fifo_in_1_5_rest_V  => fifo_in(1*NCALOFIFOS+ 5).rest,
                     fifo_in_1_6_rest_V  => fifo_in(1*NCALOFIFOS+ 6).rest,
                     fifo_in_1_7_rest_V  => fifo_in(1*NCALOFIFOS+ 7).rest,
                     fifo_in_1_8_rest_V  => fifo_in(1*NCALOFIFOS+ 8).rest,
                     fifo_in_1_9_rest_V  => fifo_in(1*NCALOFIFOS+ 9).rest,
                     fifo_in_1_10_rest_V => fifo_in(1*NCALOFIFOS+10).rest,
                     fifo_in_1_11_rest_V => fifo_in(1*NCALOFIFOS+11).rest,
                     fifo_in_1_12_rest_V => fifo_in(1*NCALOFIFOS+12).rest,
                     fifo_in_1_13_rest_V => fifo_in(1*NCALOFIFOS+13).rest,
                     fifo_in_1_14_rest_V => fifo_in(1*NCALOFIFOS+14).rest,
                     fifo_in_1_15_rest_V => fifo_in(1*NCALOFIFOS+15).rest,
                     fifo_in_1_16_rest_V => fifo_in(1*NCALOFIFOS+16).rest,
                     fifo_in_1_17_rest_V => fifo_in(1*NCALOFIFOS+17).rest,
                     fifo_in_1_18_rest_V => fifo_in(1*NCALOFIFOS+18).rest,
                     fifo_in_1_19_rest_V => fifo_in(1*NCALOFIFOS+19).rest,
                     fifo_in_2_0_rest_V  => fifo_in(2*NCALOFIFOS+ 0).rest,
                     fifo_in_2_1_rest_V  => fifo_in(2*NCALOFIFOS+ 1).rest,
                     fifo_in_2_2_rest_V  => fifo_in(2*NCALOFIFOS+ 2).rest,
                     fifo_in_2_3_rest_V  => fifo_in(2*NCALOFIFOS+ 3).rest,
                     fifo_in_2_4_rest_V  => fifo_in(2*NCALOFIFOS+ 4).rest,
                     fifo_in_2_5_rest_V  => fifo_in(2*NCALOFIFOS+ 5).rest,
                     fifo_in_2_6_rest_V  => fifo_in(2*NCALOFIFOS+ 6).rest,
                     fifo_in_2_7_rest_V  => fifo_in(2*NCALOFIFOS+ 7).rest,
                     fifo_in_2_8_rest_V  => fifo_in(2*NCALOFIFOS+ 8).rest,
                     fifo_in_2_9_rest_V  => fifo_in(2*NCALOFIFOS+ 9).rest,
                     fifo_in_2_10_rest_V => fifo_in(2*NCALOFIFOS+10).rest,
                     fifo_in_2_11_rest_V => fifo_in(2*NCALOFIFOS+11).rest,
                     fifo_in_2_12_rest_V => fifo_in(2*NCALOFIFOS+12).rest,
                     fifo_in_2_13_rest_V => fifo_in(2*NCALOFIFOS+13).rest,
                     fifo_in_2_14_rest_V => fifo_in(2*NCALOFIFOS+14).rest,
                     fifo_in_2_15_rest_V => fifo_in(2*NCALOFIFOS+15).rest,
                     fifo_in_2_16_rest_V => fifo_in(2*NCALOFIFOS+16).rest,
                     fifo_in_2_17_rest_V => fifo_in(2*NCALOFIFOS+17).rest,
                     fifo_in_2_18_rest_V => fifo_in(2*NCALOFIFOS+18).rest,
                     fifo_in_2_19_rest_V => fifo_in(2*NCALOFIFOS+19).rest,
                     fifo_out_0_0_pt_V  => fifo_out(0*NCALOFIFOS+ 0).pt,
                     fifo_out_0_1_pt_V  => fifo_out(0*NCALOFIFOS+ 1).pt,
                     fifo_out_0_2_pt_V  => fifo_out(0*NCALOFIFOS+ 2).pt,
                     fifo_out_0_3_pt_V  => fifo_out(0*NCALOFIFOS+ 3).pt,
                     fifo_out_0_4_pt_V  => fifo_out(0*NCALOFIFOS+ 4).pt,
                     fifo_out_0_5_pt_V  => fifo_out(0*NCALOFIFOS+ 5).pt,
                     fifo_out_0_6_pt_V  => fifo_out(0*NCALOFIFOS+ 6).pt,
                     fifo_out_0_7_pt_V  => fifo_out(0*NCALOFIFOS+ 7).pt,
                     fifo_out_0_8_pt_V  => fifo_out(0*NCALOFIFOS+ 8).pt,
                     fifo_out_0_9_pt_V  => fifo_out(0*NCALOFIFOS+ 9).pt,
                     fifo_out_0_10_pt_V => fifo_out(0*NCALOFIFOS+10).pt,
                     fifo_out_0_11_pt_V => fifo_out(0*NCALOFIFOS+11).pt,
                     fifo_out_0_12_pt_V => fifo_out(0*NCALOFIFOS+12).pt,
                     fifo_out_0_13_pt_V => fifo_out(0*NCALOFIFOS+13).pt,
                     fifo_out_0_14_pt_V => fifo_out(0*NCALOFIFOS+14).pt,
                     fifo_out_0_15_pt_V => fifo_out(0*NCALOFIFOS+15).pt,
                     fifo_out_0_16_pt_V => fifo_out(0*NCALOFIFOS+16).pt,
                     fifo_out_0_17_pt_V => fifo_out(0*NCALOFIFOS+17).pt,
                     fifo_out_0_18_pt_V => fifo_out(0*NCALOFIFOS+18).pt,
                     fifo_out_0_19_pt_V => fifo_out(0*NCALOFIFOS+19).pt,
                     fifo_out_1_0_pt_V  => fifo_out(1*NCALOFIFOS+ 0).pt,
                     fifo_out_1_1_pt_V  => fifo_out(1*NCALOFIFOS+ 1).pt,
                     fifo_out_1_2_pt_V  => fifo_out(1*NCALOFIFOS+ 2).pt,
                     fifo_out_1_3_pt_V  => fifo_out(1*NCALOFIFOS+ 3).pt,
                     fifo_out_1_4_pt_V  => fifo_out(1*NCALOFIFOS+ 4).pt,
                     fifo_out_1_5_pt_V  => fifo_out(1*NCALOFIFOS+ 5).pt,
                     fifo_out_1_6_pt_V  => fifo_out(1*NCALOFIFOS+ 6).pt,
                     fifo_out_1_7_pt_V  => fifo_out(1*NCALOFIFOS+ 7).pt,
                     fifo_out_1_8_pt_V  => fifo_out(1*NCALOFIFOS+ 8).pt,
                     fifo_out_1_9_pt_V  => fifo_out(1*NCALOFIFOS+ 9).pt,
                     fifo_out_1_10_pt_V => fifo_out(1*NCALOFIFOS+10).pt,
                     fifo_out_1_11_pt_V => fifo_out(1*NCALOFIFOS+11).pt,
                     fifo_out_1_12_pt_V => fifo_out(1*NCALOFIFOS+12).pt,
                     fifo_out_1_13_pt_V => fifo_out(1*NCALOFIFOS+13).pt,
                     fifo_out_1_14_pt_V => fifo_out(1*NCALOFIFOS+14).pt,
                     fifo_out_1_15_pt_V => fifo_out(1*NCALOFIFOS+15).pt,
                     fifo_out_1_16_pt_V => fifo_out(1*NCALOFIFOS+16).pt,
                     fifo_out_1_17_pt_V => fifo_out(1*NCALOFIFOS+17).pt,
                     fifo_out_1_18_pt_V => fifo_out(1*NCALOFIFOS+18).pt,
                     fifo_out_1_19_pt_V => fifo_out(1*NCALOFIFOS+19).pt,
                     fifo_out_2_0_pt_V  => fifo_out(2*NCALOFIFOS+ 0).pt,
                     fifo_out_2_1_pt_V  => fifo_out(2*NCALOFIFOS+ 1).pt,
                     fifo_out_2_2_pt_V  => fifo_out(2*NCALOFIFOS+ 2).pt,
                     fifo_out_2_3_pt_V  => fifo_out(2*NCALOFIFOS+ 3).pt,
                     fifo_out_2_4_pt_V  => fifo_out(2*NCALOFIFOS+ 4).pt,
                     fifo_out_2_5_pt_V  => fifo_out(2*NCALOFIFOS+ 5).pt,
                     fifo_out_2_6_pt_V  => fifo_out(2*NCALOFIFOS+ 6).pt,
                     fifo_out_2_7_pt_V  => fifo_out(2*NCALOFIFOS+ 7).pt,
                     fifo_out_2_8_pt_V  => fifo_out(2*NCALOFIFOS+ 8).pt,
                     fifo_out_2_9_pt_V  => fifo_out(2*NCALOFIFOS+ 9).pt,
                     fifo_out_2_10_pt_V => fifo_out(2*NCALOFIFOS+10).pt,
                     fifo_out_2_11_pt_V => fifo_out(2*NCALOFIFOS+11).pt,
                     fifo_out_2_12_pt_V => fifo_out(2*NCALOFIFOS+12).pt,
                     fifo_out_2_13_pt_V => fifo_out(2*NCALOFIFOS+13).pt,
                     fifo_out_2_14_pt_V => fifo_out(2*NCALOFIFOS+14).pt,
                     fifo_out_2_15_pt_V => fifo_out(2*NCALOFIFOS+15).pt,
                     fifo_out_2_16_pt_V => fifo_out(2*NCALOFIFOS+16).pt,
                     fifo_out_2_17_pt_V => fifo_out(2*NCALOFIFOS+17).pt,
                     fifo_out_2_18_pt_V => fifo_out(2*NCALOFIFOS+18).pt,
                     fifo_out_2_19_pt_V => fifo_out(2*NCALOFIFOS+19).pt,
                     fifo_out_0_0_eta_V  => fifo_out(0*NCALOFIFOS+ 0).eta,
                     fifo_out_0_1_eta_V  => fifo_out(0*NCALOFIFOS+ 1).eta,
                     fifo_out_0_2_eta_V  => fifo_out(0*NCALOFIFOS+ 2).eta,
                     fifo_out_0_3_eta_V  => fifo_out(0*NCALOFIFOS+ 3).eta,
                     fifo_out_0_4_eta_V  => fifo_out(0*NCALOFIFOS+ 4).eta,
                     fifo_out_0_5_eta_V  => fifo_out(0*NCALOFIFOS+ 5).eta,
                     fifo_out_0_6_eta_V  => fifo_out(0*NCALOFIFOS+ 6).eta,
                     fifo_out_0_7_eta_V  => fifo_out(0*NCALOFIFOS+ 7).eta,
                     fifo_out_0_8_eta_V  => fifo_out(0*NCALOFIFOS+ 8).eta,
                     fifo_out_0_9_eta_V  => fifo_out(0*NCALOFIFOS+ 9).eta,
                     fifo_out_0_10_eta_V => fifo_out(0*NCALOFIFOS+10).eta,
                     fifo_out_0_11_eta_V => fifo_out(0*NCALOFIFOS+11).eta,
                     fifo_out_0_12_eta_V => fifo_out(0*NCALOFIFOS+12).eta,
                     fifo_out_0_13_eta_V => fifo_out(0*NCALOFIFOS+13).eta,
                     fifo_out_0_14_eta_V => fifo_out(0*NCALOFIFOS+14).eta,
                     fifo_out_0_15_eta_V => fifo_out(0*NCALOFIFOS+15).eta,
                     fifo_out_0_16_eta_V => fifo_out(0*NCALOFIFOS+16).eta,
                     fifo_out_0_17_eta_V => fifo_out(0*NCALOFIFOS+17).eta,
                     fifo_out_0_18_eta_V => fifo_out(0*NCALOFIFOS+18).eta,
                     fifo_out_0_19_eta_V => fifo_out(0*NCALOFIFOS+19).eta,
                     fifo_out_1_0_eta_V  => fifo_out(1*NCALOFIFOS+ 0).eta,
                     fifo_out_1_1_eta_V  => fifo_out(1*NCALOFIFOS+ 1).eta,
                     fifo_out_1_2_eta_V  => fifo_out(1*NCALOFIFOS+ 2).eta,
                     fifo_out_1_3_eta_V  => fifo_out(1*NCALOFIFOS+ 3).eta,
                     fifo_out_1_4_eta_V  => fifo_out(1*NCALOFIFOS+ 4).eta,
                     fifo_out_1_5_eta_V  => fifo_out(1*NCALOFIFOS+ 5).eta,
                     fifo_out_1_6_eta_V  => fifo_out(1*NCALOFIFOS+ 6).eta,
                     fifo_out_1_7_eta_V  => fifo_out(1*NCALOFIFOS+ 7).eta,
                     fifo_out_1_8_eta_V  => fifo_out(1*NCALOFIFOS+ 8).eta,
                     fifo_out_1_9_eta_V  => fifo_out(1*NCALOFIFOS+ 9).eta,
                     fifo_out_1_10_eta_V => fifo_out(1*NCALOFIFOS+10).eta,
                     fifo_out_1_11_eta_V => fifo_out(1*NCALOFIFOS+11).eta,
                     fifo_out_1_12_eta_V => fifo_out(1*NCALOFIFOS+12).eta,
                     fifo_out_1_13_eta_V => fifo_out(1*NCALOFIFOS+13).eta,
                     fifo_out_1_14_eta_V => fifo_out(1*NCALOFIFOS+14).eta,
                     fifo_out_1_15_eta_V => fifo_out(1*NCALOFIFOS+15).eta,
                     fifo_out_1_16_eta_V => fifo_out(1*NCALOFIFOS+16).eta,
                     fifo_out_1_17_eta_V => fifo_out(1*NCALOFIFOS+17).eta,
                     fifo_out_1_18_eta_V => fifo_out(1*NCALOFIFOS+18).eta,
                     fifo_out_1_19_eta_V => fifo_out(1*NCALOFIFOS+19).eta,
                     fifo_out_2_0_eta_V  => fifo_out(2*NCALOFIFOS+ 0).eta,
                     fifo_out_2_1_eta_V  => fifo_out(2*NCALOFIFOS+ 1).eta,
                     fifo_out_2_2_eta_V  => fifo_out(2*NCALOFIFOS+ 2).eta,
                     fifo_out_2_3_eta_V  => fifo_out(2*NCALOFIFOS+ 3).eta,
                     fifo_out_2_4_eta_V  => fifo_out(2*NCALOFIFOS+ 4).eta,
                     fifo_out_2_5_eta_V  => fifo_out(2*NCALOFIFOS+ 5).eta,
                     fifo_out_2_6_eta_V  => fifo_out(2*NCALOFIFOS+ 6).eta,
                     fifo_out_2_7_eta_V  => fifo_out(2*NCALOFIFOS+ 7).eta,
                     fifo_out_2_8_eta_V  => fifo_out(2*NCALOFIFOS+ 8).eta,
                     fifo_out_2_9_eta_V  => fifo_out(2*NCALOFIFOS+ 9).eta,
                     fifo_out_2_10_eta_V => fifo_out(2*NCALOFIFOS+10).eta,
                     fifo_out_2_11_eta_V => fifo_out(2*NCALOFIFOS+11).eta,
                     fifo_out_2_12_eta_V => fifo_out(2*NCALOFIFOS+12).eta,
                     fifo_out_2_13_eta_V => fifo_out(2*NCALOFIFOS+13).eta,
                     fifo_out_2_14_eta_V => fifo_out(2*NCALOFIFOS+14).eta,
                     fifo_out_2_15_eta_V => fifo_out(2*NCALOFIFOS+15).eta,
                     fifo_out_2_16_eta_V => fifo_out(2*NCALOFIFOS+16).eta,
                     fifo_out_2_17_eta_V => fifo_out(2*NCALOFIFOS+17).eta,
                     fifo_out_2_18_eta_V => fifo_out(2*NCALOFIFOS+18).eta,
                     fifo_out_2_19_eta_V => fifo_out(2*NCALOFIFOS+19).eta,
                     fifo_out_0_0_phi_V  => fifo_out(0*NCALOFIFOS+ 0).phi,
                     fifo_out_0_1_phi_V  => fifo_out(0*NCALOFIFOS+ 1).phi,
                     fifo_out_0_2_phi_V  => fifo_out(0*NCALOFIFOS+ 2).phi,
                     fifo_out_0_3_phi_V  => fifo_out(0*NCALOFIFOS+ 3).phi,
                     fifo_out_0_4_phi_V  => fifo_out(0*NCALOFIFOS+ 4).phi,
                     fifo_out_0_5_phi_V  => fifo_out(0*NCALOFIFOS+ 5).phi,
                     fifo_out_0_6_phi_V  => fifo_out(0*NCALOFIFOS+ 6).phi,
                     fifo_out_0_7_phi_V  => fifo_out(0*NCALOFIFOS+ 7).phi,
                     fifo_out_0_8_phi_V  => fifo_out(0*NCALOFIFOS+ 8).phi,
                     fifo_out_0_9_phi_V  => fifo_out(0*NCALOFIFOS+ 9).phi,
                     fifo_out_0_10_phi_V => fifo_out(0*NCALOFIFOS+10).phi,
                     fifo_out_0_11_phi_V => fifo_out(0*NCALOFIFOS+11).phi,
                     fifo_out_0_12_phi_V => fifo_out(0*NCALOFIFOS+12).phi,
                     fifo_out_0_13_phi_V => fifo_out(0*NCALOFIFOS+13).phi,
                     fifo_out_0_14_phi_V => fifo_out(0*NCALOFIFOS+14).phi,
                     fifo_out_0_15_phi_V => fifo_out(0*NCALOFIFOS+15).phi,
                     fifo_out_0_16_phi_V => fifo_out(0*NCALOFIFOS+16).phi,
                     fifo_out_0_17_phi_V => fifo_out(0*NCALOFIFOS+17).phi,
                     fifo_out_0_18_phi_V => fifo_out(0*NCALOFIFOS+18).phi,
                     fifo_out_0_19_phi_V => fifo_out(0*NCALOFIFOS+19).phi,
                     fifo_out_1_0_phi_V  => fifo_out(1*NCALOFIFOS+ 0).phi,
                     fifo_out_1_1_phi_V  => fifo_out(1*NCALOFIFOS+ 1).phi,
                     fifo_out_1_2_phi_V  => fifo_out(1*NCALOFIFOS+ 2).phi,
                     fifo_out_1_3_phi_V  => fifo_out(1*NCALOFIFOS+ 3).phi,
                     fifo_out_1_4_phi_V  => fifo_out(1*NCALOFIFOS+ 4).phi,
                     fifo_out_1_5_phi_V  => fifo_out(1*NCALOFIFOS+ 5).phi,
                     fifo_out_1_6_phi_V  => fifo_out(1*NCALOFIFOS+ 6).phi,
                     fifo_out_1_7_phi_V  => fifo_out(1*NCALOFIFOS+ 7).phi,
                     fifo_out_1_8_phi_V  => fifo_out(1*NCALOFIFOS+ 8).phi,
                     fifo_out_1_9_phi_V  => fifo_out(1*NCALOFIFOS+ 9).phi,
                     fifo_out_1_10_phi_V => fifo_out(1*NCALOFIFOS+10).phi,
                     fifo_out_1_11_phi_V => fifo_out(1*NCALOFIFOS+11).phi,
                     fifo_out_1_12_phi_V => fifo_out(1*NCALOFIFOS+12).phi,
                     fifo_out_1_13_phi_V => fifo_out(1*NCALOFIFOS+13).phi,
                     fifo_out_1_14_phi_V => fifo_out(1*NCALOFIFOS+14).phi,
                     fifo_out_1_15_phi_V => fifo_out(1*NCALOFIFOS+15).phi,
                     fifo_out_1_16_phi_V => fifo_out(1*NCALOFIFOS+16).phi,
                     fifo_out_1_17_phi_V => fifo_out(1*NCALOFIFOS+17).phi,
                     fifo_out_1_18_phi_V => fifo_out(1*NCALOFIFOS+18).phi,
                     fifo_out_1_19_phi_V => fifo_out(1*NCALOFIFOS+19).phi,
                     fifo_out_2_0_phi_V  => fifo_out(2*NCALOFIFOS+ 0).phi,
                     fifo_out_2_1_phi_V  => fifo_out(2*NCALOFIFOS+ 1).phi,
                     fifo_out_2_2_phi_V  => fifo_out(2*NCALOFIFOS+ 2).phi,
                     fifo_out_2_3_phi_V  => fifo_out(2*NCALOFIFOS+ 3).phi,
                     fifo_out_2_4_phi_V  => fifo_out(2*NCALOFIFOS+ 4).phi,
                     fifo_out_2_5_phi_V  => fifo_out(2*NCALOFIFOS+ 5).phi,
                     fifo_out_2_6_phi_V  => fifo_out(2*NCALOFIFOS+ 6).phi,
                     fifo_out_2_7_phi_V  => fifo_out(2*NCALOFIFOS+ 7).phi,
                     fifo_out_2_8_phi_V  => fifo_out(2*NCALOFIFOS+ 8).phi,
                     fifo_out_2_9_phi_V  => fifo_out(2*NCALOFIFOS+ 9).phi,
                     fifo_out_2_10_phi_V => fifo_out(2*NCALOFIFOS+10).phi,
                     fifo_out_2_11_phi_V => fifo_out(2*NCALOFIFOS+11).phi,
                     fifo_out_2_12_phi_V => fifo_out(2*NCALOFIFOS+12).phi,
                     fifo_out_2_13_phi_V => fifo_out(2*NCALOFIFOS+13).phi,
                     fifo_out_2_14_phi_V => fifo_out(2*NCALOFIFOS+14).phi,
                     fifo_out_2_15_phi_V => fifo_out(2*NCALOFIFOS+15).phi,
                     fifo_out_2_16_phi_V => fifo_out(2*NCALOFIFOS+16).phi,
                     fifo_out_2_17_phi_V => fifo_out(2*NCALOFIFOS+17).phi,
                     fifo_out_2_18_phi_V => fifo_out(2*NCALOFIFOS+18).phi,
                     fifo_out_2_19_phi_V => fifo_out(2*NCALOFIFOS+19).phi,
                     fifo_out_0_0_rest_V  => fifo_out(0*NCALOFIFOS+ 0).rest,
                     fifo_out_0_1_rest_V  => fifo_out(0*NCALOFIFOS+ 1).rest,
                     fifo_out_0_2_rest_V  => fifo_out(0*NCALOFIFOS+ 2).rest,
                     fifo_out_0_3_rest_V  => fifo_out(0*NCALOFIFOS+ 3).rest,
                     fifo_out_0_4_rest_V  => fifo_out(0*NCALOFIFOS+ 4).rest,
                     fifo_out_0_5_rest_V  => fifo_out(0*NCALOFIFOS+ 5).rest,
                     fifo_out_0_6_rest_V  => fifo_out(0*NCALOFIFOS+ 6).rest,
                     fifo_out_0_7_rest_V  => fifo_out(0*NCALOFIFOS+ 7).rest,
                     fifo_out_0_8_rest_V  => fifo_out(0*NCALOFIFOS+ 8).rest,
                     fifo_out_0_9_rest_V  => fifo_out(0*NCALOFIFOS+ 9).rest,
                     fifo_out_0_10_rest_V => fifo_out(0*NCALOFIFOS+10).rest,
                     fifo_out_0_11_rest_V => fifo_out(0*NCALOFIFOS+11).rest,
                     fifo_out_0_12_rest_V => fifo_out(0*NCALOFIFOS+12).rest,
                     fifo_out_0_13_rest_V => fifo_out(0*NCALOFIFOS+13).rest,
                     fifo_out_0_14_rest_V => fifo_out(0*NCALOFIFOS+14).rest,
                     fifo_out_0_15_rest_V => fifo_out(0*NCALOFIFOS+15).rest,
                     fifo_out_0_16_rest_V => fifo_out(0*NCALOFIFOS+16).rest,
                     fifo_out_0_17_rest_V => fifo_out(0*NCALOFIFOS+17).rest,
                     fifo_out_0_18_rest_V => fifo_out(0*NCALOFIFOS+18).rest,
                     fifo_out_0_19_rest_V => fifo_out(0*NCALOFIFOS+19).rest,
                     fifo_out_1_0_rest_V  => fifo_out(1*NCALOFIFOS+ 0).rest,
                     fifo_out_1_1_rest_V  => fifo_out(1*NCALOFIFOS+ 1).rest,
                     fifo_out_1_2_rest_V  => fifo_out(1*NCALOFIFOS+ 2).rest,
                     fifo_out_1_3_rest_V  => fifo_out(1*NCALOFIFOS+ 3).rest,
                     fifo_out_1_4_rest_V  => fifo_out(1*NCALOFIFOS+ 4).rest,
                     fifo_out_1_5_rest_V  => fifo_out(1*NCALOFIFOS+ 5).rest,
                     fifo_out_1_6_rest_V  => fifo_out(1*NCALOFIFOS+ 6).rest,
                     fifo_out_1_7_rest_V  => fifo_out(1*NCALOFIFOS+ 7).rest,
                     fifo_out_1_8_rest_V  => fifo_out(1*NCALOFIFOS+ 8).rest,
                     fifo_out_1_9_rest_V  => fifo_out(1*NCALOFIFOS+ 9).rest,
                     fifo_out_1_10_rest_V => fifo_out(1*NCALOFIFOS+10).rest,
                     fifo_out_1_11_rest_V => fifo_out(1*NCALOFIFOS+11).rest,
                     fifo_out_1_12_rest_V => fifo_out(1*NCALOFIFOS+12).rest,
                     fifo_out_1_13_rest_V => fifo_out(1*NCALOFIFOS+13).rest,
                     fifo_out_1_14_rest_V => fifo_out(1*NCALOFIFOS+14).rest,
                     fifo_out_1_15_rest_V => fifo_out(1*NCALOFIFOS+15).rest,
                     fifo_out_1_16_rest_V => fifo_out(1*NCALOFIFOS+16).rest,
                     fifo_out_1_17_rest_V => fifo_out(1*NCALOFIFOS+17).rest,
                     fifo_out_1_18_rest_V => fifo_out(1*NCALOFIFOS+18).rest,
                     fifo_out_1_19_rest_V => fifo_out(1*NCALOFIFOS+19).rest,
                     fifo_out_2_0_rest_V  => fifo_out(2*NCALOFIFOS+ 0).rest,
                     fifo_out_2_1_rest_V  => fifo_out(2*NCALOFIFOS+ 1).rest,
                     fifo_out_2_2_rest_V  => fifo_out(2*NCALOFIFOS+ 2).rest,
                     fifo_out_2_3_rest_V  => fifo_out(2*NCALOFIFOS+ 3).rest,
                     fifo_out_2_4_rest_V  => fifo_out(2*NCALOFIFOS+ 4).rest,
                     fifo_out_2_5_rest_V  => fifo_out(2*NCALOFIFOS+ 5).rest,
                     fifo_out_2_6_rest_V  => fifo_out(2*NCALOFIFOS+ 6).rest,
                     fifo_out_2_7_rest_V  => fifo_out(2*NCALOFIFOS+ 7).rest,
                     fifo_out_2_8_rest_V  => fifo_out(2*NCALOFIFOS+ 8).rest,
                     fifo_out_2_9_rest_V  => fifo_out(2*NCALOFIFOS+ 9).rest,
                     fifo_out_2_10_rest_V => fifo_out(2*NCALOFIFOS+10).rest,
                     fifo_out_2_11_rest_V => fifo_out(2*NCALOFIFOS+11).rest,
                     fifo_out_2_12_rest_V => fifo_out(2*NCALOFIFOS+12).rest,
                     fifo_out_2_13_rest_V => fifo_out(2*NCALOFIFOS+13).rest,
                     fifo_out_2_14_rest_V => fifo_out(2*NCALOFIFOS+14).rest,
                     fifo_out_2_15_rest_V => fifo_out(2*NCALOFIFOS+15).rest,
                     fifo_out_2_16_rest_V => fifo_out(2*NCALOFIFOS+16).rest,
                     fifo_out_2_17_rest_V => fifo_out(2*NCALOFIFOS+17).rest,
                     fifo_out_2_18_rest_V => fifo_out(2*NCALOFIFOS+18).rest,
                     fifo_out_2_19_rest_V => fifo_out(2*NCALOFIFOS+19).rest,
                     fifo_write_0_0  => fifo_write(0*NCALOFIFOS+ 0),
                     fifo_write_0_1  => fifo_write(0*NCALOFIFOS+ 1),
                     fifo_write_0_2  => fifo_write(0*NCALOFIFOS+ 2),
                     fifo_write_0_3  => fifo_write(0*NCALOFIFOS+ 3),
                     fifo_write_0_4  => fifo_write(0*NCALOFIFOS+ 4),
                     fifo_write_0_5  => fifo_write(0*NCALOFIFOS+ 5),
                     fifo_write_0_6  => fifo_write(0*NCALOFIFOS+ 6),
                     fifo_write_0_7  => fifo_write(0*NCALOFIFOS+ 7),
                     fifo_write_0_8  => fifo_write(0*NCALOFIFOS+ 8),
                     fifo_write_0_9  => fifo_write(0*NCALOFIFOS+ 9),
                     fifo_write_0_10 => fifo_write(0*NCALOFIFOS+10),
                     fifo_write_0_11 => fifo_write(0*NCALOFIFOS+11),
                     fifo_write_0_12 => fifo_write(0*NCALOFIFOS+12),
                     fifo_write_0_13 => fifo_write(0*NCALOFIFOS+13),
                     fifo_write_0_14 => fifo_write(0*NCALOFIFOS+14),
                     fifo_write_0_15 => fifo_write(0*NCALOFIFOS+15),
                     fifo_write_0_16 => fifo_write(0*NCALOFIFOS+16),
                     fifo_write_0_17 => fifo_write(0*NCALOFIFOS+17),
                     fifo_write_0_18 => fifo_write(0*NCALOFIFOS+18),
                     fifo_write_0_19 => fifo_write(0*NCALOFIFOS+19),
                     fifo_write_1_0  => fifo_write(1*NCALOFIFOS+ 0),
                     fifo_write_1_1  => fifo_write(1*NCALOFIFOS+ 1),
                     fifo_write_1_2  => fifo_write(1*NCALOFIFOS+ 2),
                     fifo_write_1_3  => fifo_write(1*NCALOFIFOS+ 3),
                     fifo_write_1_4  => fifo_write(1*NCALOFIFOS+ 4),
                     fifo_write_1_5  => fifo_write(1*NCALOFIFOS+ 5),
                     fifo_write_1_6  => fifo_write(1*NCALOFIFOS+ 6),
                     fifo_write_1_7  => fifo_write(1*NCALOFIFOS+ 7),
                     fifo_write_1_8  => fifo_write(1*NCALOFIFOS+ 8),
                     fifo_write_1_9  => fifo_write(1*NCALOFIFOS+ 9),
                     fifo_write_1_10 => fifo_write(1*NCALOFIFOS+10),
                     fifo_write_1_11 => fifo_write(1*NCALOFIFOS+11),
                     fifo_write_1_12 => fifo_write(1*NCALOFIFOS+12),
                     fifo_write_1_13 => fifo_write(1*NCALOFIFOS+13),
                     fifo_write_1_14 => fifo_write(1*NCALOFIFOS+14),
                     fifo_write_1_15 => fifo_write(1*NCALOFIFOS+15),
                     fifo_write_1_16 => fifo_write(1*NCALOFIFOS+16),
                     fifo_write_1_17 => fifo_write(1*NCALOFIFOS+17),
                     fifo_write_1_18 => fifo_write(1*NCALOFIFOS+18),
                     fifo_write_1_19 => fifo_write(1*NCALOFIFOS+19),
                     fifo_write_2_0  => fifo_write(2*NCALOFIFOS+ 0),
                     fifo_write_2_1  => fifo_write(2*NCALOFIFOS+ 1),
                     fifo_write_2_2  => fifo_write(2*NCALOFIFOS+ 2),
                     fifo_write_2_3  => fifo_write(2*NCALOFIFOS+ 3),
                     fifo_write_2_4  => fifo_write(2*NCALOFIFOS+ 4),
                     fifo_write_2_5  => fifo_write(2*NCALOFIFOS+ 5),
                     fifo_write_2_6  => fifo_write(2*NCALOFIFOS+ 6),
                     fifo_write_2_7  => fifo_write(2*NCALOFIFOS+ 7),
                     fifo_write_2_8  => fifo_write(2*NCALOFIFOS+ 8),
                     fifo_write_2_9  => fifo_write(2*NCALOFIFOS+ 9),
                     fifo_write_2_10 => fifo_write(2*NCALOFIFOS+10),
                     fifo_write_2_11 => fifo_write(2*NCALOFIFOS+11),
                     fifo_write_2_12 => fifo_write(2*NCALOFIFOS+12),
                     fifo_write_2_13 => fifo_write(2*NCALOFIFOS+13),
                     fifo_write_2_14 => fifo_write(2*NCALOFIFOS+14),
                     fifo_write_2_15 => fifo_write(2*NCALOFIFOS+15),
                     fifo_write_2_16 => fifo_write(2*NCALOFIFOS+16),
                     fifo_write_2_17 => fifo_write(2*NCALOFIFOS+17),
                     fifo_write_2_18 => fifo_write(2*NCALOFIFOS+18),
                     fifo_write_2_19 => fifo_write(2*NCALOFIFOS+19),
                     fifo_full_0_0  => fifo_full(0*NCALOFIFOS+ 0),
                     fifo_full_0_1  => fifo_full(0*NCALOFIFOS+ 1),
                     fifo_full_0_2  => fifo_full(0*NCALOFIFOS+ 2),
                     fifo_full_0_3  => fifo_full(0*NCALOFIFOS+ 3),
                     fifo_full_0_4  => fifo_full(0*NCALOFIFOS+ 4),
                     fifo_full_0_5  => fifo_full(0*NCALOFIFOS+ 5),
                     fifo_full_0_6  => fifo_full(0*NCALOFIFOS+ 6),
                     fifo_full_0_7  => fifo_full(0*NCALOFIFOS+ 7),
                     fifo_full_0_8  => fifo_full(0*NCALOFIFOS+ 8),
                     fifo_full_0_9  => fifo_full(0*NCALOFIFOS+ 9),
                     fifo_full_0_10 => fifo_full(0*NCALOFIFOS+10),
                     fifo_full_0_11 => fifo_full(0*NCALOFIFOS+11),
                     fifo_full_0_12 => fifo_full(0*NCALOFIFOS+12),
                     fifo_full_0_13 => fifo_full(0*NCALOFIFOS+13),
                     fifo_full_0_14 => fifo_full(0*NCALOFIFOS+14),
                     fifo_full_0_15 => fifo_full(0*NCALOFIFOS+15),
                     fifo_full_0_16 => fifo_full(0*NCALOFIFOS+16),
                     fifo_full_0_17 => fifo_full(0*NCALOFIFOS+17),
                     fifo_full_0_18 => fifo_full(0*NCALOFIFOS+18),
                     fifo_full_0_19 => fifo_full(0*NCALOFIFOS+19),
                     fifo_full_1_0  => fifo_full(1*NCALOFIFOS+ 0),
                     fifo_full_1_1  => fifo_full(1*NCALOFIFOS+ 1),
                     fifo_full_1_2  => fifo_full(1*NCALOFIFOS+ 2),
                     fifo_full_1_3  => fifo_full(1*NCALOFIFOS+ 3),
                     fifo_full_1_4  => fifo_full(1*NCALOFIFOS+ 4),
                     fifo_full_1_5  => fifo_full(1*NCALOFIFOS+ 5),
                     fifo_full_1_6  => fifo_full(1*NCALOFIFOS+ 6),
                     fifo_full_1_7  => fifo_full(1*NCALOFIFOS+ 7),
                     fifo_full_1_8  => fifo_full(1*NCALOFIFOS+ 8),
                     fifo_full_1_9  => fifo_full(1*NCALOFIFOS+ 9),
                     fifo_full_1_10 => fifo_full(1*NCALOFIFOS+10),
                     fifo_full_1_11 => fifo_full(1*NCALOFIFOS+11),
                     fifo_full_1_12 => fifo_full(1*NCALOFIFOS+12),
                     fifo_full_1_13 => fifo_full(1*NCALOFIFOS+13),
                     fifo_full_1_14 => fifo_full(1*NCALOFIFOS+14),
                     fifo_full_1_15 => fifo_full(1*NCALOFIFOS+15),
                     fifo_full_1_16 => fifo_full(1*NCALOFIFOS+16),
                     fifo_full_1_17 => fifo_full(1*NCALOFIFOS+17),
                     fifo_full_1_18 => fifo_full(1*NCALOFIFOS+18),
                     fifo_full_1_19 => fifo_full(1*NCALOFIFOS+19),
                     fifo_full_2_0  => fifo_full(2*NCALOFIFOS+ 0),
                     fifo_full_2_1  => fifo_full(2*NCALOFIFOS+ 1),
                     fifo_full_2_2  => fifo_full(2*NCALOFIFOS+ 2),
                     fifo_full_2_3  => fifo_full(2*NCALOFIFOS+ 3),
                     fifo_full_2_4  => fifo_full(2*NCALOFIFOS+ 4),
                     fifo_full_2_5  => fifo_full(2*NCALOFIFOS+ 5),
                     fifo_full_2_6  => fifo_full(2*NCALOFIFOS+ 6),
                     fifo_full_2_7  => fifo_full(2*NCALOFIFOS+ 7),
                     fifo_full_2_8  => fifo_full(2*NCALOFIFOS+ 8),
                     fifo_full_2_9  => fifo_full(2*NCALOFIFOS+ 9),
                     fifo_full_2_10 => fifo_full(2*NCALOFIFOS+10),
                     fifo_full_2_11 => fifo_full(2*NCALOFIFOS+11),
                     fifo_full_2_12 => fifo_full(2*NCALOFIFOS+12),
                     fifo_full_2_13 => fifo_full(2*NCALOFIFOS+13),
                     fifo_full_2_14 => fifo_full(2*NCALOFIFOS+14),
                     fifo_full_2_15 => fifo_full(2*NCALOFIFOS+15),
                     fifo_full_2_16 => fifo_full(2*NCALOFIFOS+16),
                     fifo_full_2_17 => fifo_full(2*NCALOFIFOS+17),
                     fifo_full_2_18 => fifo_full(2*NCALOFIFOS+18),
                     fifo_full_2_19 => fifo_full(2*NCALOFIFOS+19),
                     fifo_out_valid_0_0  => fifo_out_valid(0*NCALOFIFOS+ 0),
                     fifo_out_valid_0_1  => fifo_out_valid(0*NCALOFIFOS+ 1),
                     fifo_out_valid_0_2  => fifo_out_valid(0*NCALOFIFOS+ 2),
                     fifo_out_valid_0_3  => fifo_out_valid(0*NCALOFIFOS+ 3),
                     fifo_out_valid_0_4  => fifo_out_valid(0*NCALOFIFOS+ 4),
                     fifo_out_valid_0_5  => fifo_out_valid(0*NCALOFIFOS+ 5),
                     fifo_out_valid_0_6  => fifo_out_valid(0*NCALOFIFOS+ 6),
                     fifo_out_valid_0_7  => fifo_out_valid(0*NCALOFIFOS+ 7),
                     fifo_out_valid_0_8  => fifo_out_valid(0*NCALOFIFOS+ 8),
                     fifo_out_valid_0_9  => fifo_out_valid(0*NCALOFIFOS+ 9),
                     fifo_out_valid_0_10 => fifo_out_valid(0*NCALOFIFOS+10),
                     fifo_out_valid_0_11 => fifo_out_valid(0*NCALOFIFOS+11),
                     fifo_out_valid_0_12 => fifo_out_valid(0*NCALOFIFOS+12),
                     fifo_out_valid_0_13 => fifo_out_valid(0*NCALOFIFOS+13),
                     fifo_out_valid_0_14 => fifo_out_valid(0*NCALOFIFOS+14),
                     fifo_out_valid_0_15 => fifo_out_valid(0*NCALOFIFOS+15),
                     fifo_out_valid_0_16 => fifo_out_valid(0*NCALOFIFOS+16),
                     fifo_out_valid_0_17 => fifo_out_valid(0*NCALOFIFOS+17),
                     fifo_out_valid_0_18 => fifo_out_valid(0*NCALOFIFOS+18),
                     fifo_out_valid_0_19 => fifo_out_valid(0*NCALOFIFOS+19),
                     fifo_out_valid_1_0  => fifo_out_valid(1*NCALOFIFOS+ 0),
                     fifo_out_valid_1_1  => fifo_out_valid(1*NCALOFIFOS+ 1),
                     fifo_out_valid_1_2  => fifo_out_valid(1*NCALOFIFOS+ 2),
                     fifo_out_valid_1_3  => fifo_out_valid(1*NCALOFIFOS+ 3),
                     fifo_out_valid_1_4  => fifo_out_valid(1*NCALOFIFOS+ 4),
                     fifo_out_valid_1_5  => fifo_out_valid(1*NCALOFIFOS+ 5),
                     fifo_out_valid_1_6  => fifo_out_valid(1*NCALOFIFOS+ 6),
                     fifo_out_valid_1_7  => fifo_out_valid(1*NCALOFIFOS+ 7),
                     fifo_out_valid_1_8  => fifo_out_valid(1*NCALOFIFOS+ 8),
                     fifo_out_valid_1_9  => fifo_out_valid(1*NCALOFIFOS+ 9),
                     fifo_out_valid_1_10 => fifo_out_valid(1*NCALOFIFOS+10),
                     fifo_out_valid_1_11 => fifo_out_valid(1*NCALOFIFOS+11),
                     fifo_out_valid_1_12 => fifo_out_valid(1*NCALOFIFOS+12),
                     fifo_out_valid_1_13 => fifo_out_valid(1*NCALOFIFOS+13),
                     fifo_out_valid_1_14 => fifo_out_valid(1*NCALOFIFOS+14),
                     fifo_out_valid_1_15 => fifo_out_valid(1*NCALOFIFOS+15),
                     fifo_out_valid_1_16 => fifo_out_valid(1*NCALOFIFOS+16),
                     fifo_out_valid_1_17 => fifo_out_valid(1*NCALOFIFOS+17),
                     fifo_out_valid_1_18 => fifo_out_valid(1*NCALOFIFOS+18),
                     fifo_out_valid_1_19 => fifo_out_valid(1*NCALOFIFOS+19),
                     fifo_out_valid_2_0  => fifo_out_valid(2*NCALOFIFOS+ 0),
                     fifo_out_valid_2_1  => fifo_out_valid(2*NCALOFIFOS+ 1),
                     fifo_out_valid_2_2  => fifo_out_valid(2*NCALOFIFOS+ 2),
                     fifo_out_valid_2_3  => fifo_out_valid(2*NCALOFIFOS+ 3),
                     fifo_out_valid_2_4  => fifo_out_valid(2*NCALOFIFOS+ 4),
                     fifo_out_valid_2_5  => fifo_out_valid(2*NCALOFIFOS+ 5),
                     fifo_out_valid_2_6  => fifo_out_valid(2*NCALOFIFOS+ 6),
                     fifo_out_valid_2_7  => fifo_out_valid(2*NCALOFIFOS+ 7),
                     fifo_out_valid_2_8  => fifo_out_valid(2*NCALOFIFOS+ 8),
                     fifo_out_valid_2_9  => fifo_out_valid(2*NCALOFIFOS+ 9),
                     fifo_out_valid_2_10 => fifo_out_valid(2*NCALOFIFOS+10),
                     fifo_out_valid_2_11 => fifo_out_valid(2*NCALOFIFOS+11),
                     fifo_out_valid_2_12 => fifo_out_valid(2*NCALOFIFOS+12),
                     fifo_out_valid_2_13 => fifo_out_valid(2*NCALOFIFOS+13),
                     fifo_out_valid_2_14 => fifo_out_valid(2*NCALOFIFOS+14),
                     fifo_out_valid_2_15 => fifo_out_valid(2*NCALOFIFOS+15),
                     fifo_out_valid_2_16 => fifo_out_valid(2*NCALOFIFOS+16),
                     fifo_out_valid_2_17 => fifo_out_valid(2*NCALOFIFOS+17),
                     fifo_out_valid_2_18 => fifo_out_valid(2*NCALOFIFOS+18),
                     fifo_out_valid_2_19 => fifo_out_valid(2*NCALOFIFOS+19),
                     fifo_out_roll_0_0  => fifo_out_roll(0*NCALOFIFOS+ 0),
                     fifo_out_roll_0_1  => fifo_out_roll(0*NCALOFIFOS+ 1),
                     fifo_out_roll_0_2  => fifo_out_roll(0*NCALOFIFOS+ 2),
                     fifo_out_roll_0_3  => fifo_out_roll(0*NCALOFIFOS+ 3),
                     fifo_out_roll_0_4  => fifo_out_roll(0*NCALOFIFOS+ 4),
                     fifo_out_roll_0_5  => fifo_out_roll(0*NCALOFIFOS+ 5),
                     fifo_out_roll_0_6  => fifo_out_roll(0*NCALOFIFOS+ 6),
                     fifo_out_roll_0_7  => fifo_out_roll(0*NCALOFIFOS+ 7),
                     fifo_out_roll_0_8  => fifo_out_roll(0*NCALOFIFOS+ 8),
                     fifo_out_roll_0_9  => fifo_out_roll(0*NCALOFIFOS+ 9),
                     fifo_out_roll_0_10 => fifo_out_roll(0*NCALOFIFOS+10),
                     fifo_out_roll_0_11 => fifo_out_roll(0*NCALOFIFOS+11),
                     fifo_out_roll_0_12 => fifo_out_roll(0*NCALOFIFOS+12),
                     fifo_out_roll_0_13 => fifo_out_roll(0*NCALOFIFOS+13),
                     fifo_out_roll_0_14 => fifo_out_roll(0*NCALOFIFOS+14),
                     fifo_out_roll_0_15 => fifo_out_roll(0*NCALOFIFOS+15),
                     fifo_out_roll_0_16 => fifo_out_roll(0*NCALOFIFOS+16),
                     fifo_out_roll_0_17 => fifo_out_roll(0*NCALOFIFOS+17),
                     fifo_out_roll_0_18 => fifo_out_roll(0*NCALOFIFOS+18),
                     fifo_out_roll_0_19 => fifo_out_roll(0*NCALOFIFOS+19),
                     fifo_out_roll_1_0  => fifo_out_roll(1*NCALOFIFOS+ 0),
                     fifo_out_roll_1_1  => fifo_out_roll(1*NCALOFIFOS+ 1),
                     fifo_out_roll_1_2  => fifo_out_roll(1*NCALOFIFOS+ 2),
                     fifo_out_roll_1_3  => fifo_out_roll(1*NCALOFIFOS+ 3),
                     fifo_out_roll_1_4  => fifo_out_roll(1*NCALOFIFOS+ 4),
                     fifo_out_roll_1_5  => fifo_out_roll(1*NCALOFIFOS+ 5),
                     fifo_out_roll_1_6  => fifo_out_roll(1*NCALOFIFOS+ 6),
                     fifo_out_roll_1_7  => fifo_out_roll(1*NCALOFIFOS+ 7),
                     fifo_out_roll_1_8  => fifo_out_roll(1*NCALOFIFOS+ 8),
                     fifo_out_roll_1_9  => fifo_out_roll(1*NCALOFIFOS+ 9),
                     fifo_out_roll_1_10 => fifo_out_roll(1*NCALOFIFOS+10),
                     fifo_out_roll_1_11 => fifo_out_roll(1*NCALOFIFOS+11),
                     fifo_out_roll_1_12 => fifo_out_roll(1*NCALOFIFOS+12),
                     fifo_out_roll_1_13 => fifo_out_roll(1*NCALOFIFOS+13),
                     fifo_out_roll_1_14 => fifo_out_roll(1*NCALOFIFOS+14),
                     fifo_out_roll_1_15 => fifo_out_roll(1*NCALOFIFOS+15),
                     fifo_out_roll_1_16 => fifo_out_roll(1*NCALOFIFOS+16),
                     fifo_out_roll_1_17 => fifo_out_roll(1*NCALOFIFOS+17),
                     fifo_out_roll_1_18 => fifo_out_roll(1*NCALOFIFOS+18),
                     fifo_out_roll_1_19 => fifo_out_roll(1*NCALOFIFOS+19),
                     fifo_out_roll_2_0  => fifo_out_roll(2*NCALOFIFOS+ 0),
                     fifo_out_roll_2_1  => fifo_out_roll(2*NCALOFIFOS+ 1),
                     fifo_out_roll_2_2  => fifo_out_roll(2*NCALOFIFOS+ 2),
                     fifo_out_roll_2_3  => fifo_out_roll(2*NCALOFIFOS+ 3),
                     fifo_out_roll_2_4  => fifo_out_roll(2*NCALOFIFOS+ 4),
                     fifo_out_roll_2_5  => fifo_out_roll(2*NCALOFIFOS+ 5),
                     fifo_out_roll_2_6  => fifo_out_roll(2*NCALOFIFOS+ 6),
                     fifo_out_roll_2_7  => fifo_out_roll(2*NCALOFIFOS+ 7),
                     fifo_out_roll_2_8  => fifo_out_roll(2*NCALOFIFOS+ 8),
                     fifo_out_roll_2_9  => fifo_out_roll(2*NCALOFIFOS+ 9),
                     fifo_out_roll_2_10 => fifo_out_roll(2*NCALOFIFOS+10),
                     fifo_out_roll_2_11 => fifo_out_roll(2*NCALOFIFOS+11),
                     fifo_out_roll_2_12 => fifo_out_roll(2*NCALOFIFOS+12),
                     fifo_out_roll_2_13 => fifo_out_roll(2*NCALOFIFOS+13),
                     fifo_out_roll_2_14 => fifo_out_roll(2*NCALOFIFOS+14),
                     fifo_out_roll_2_15 => fifo_out_roll(2*NCALOFIFOS+15),
                     fifo_out_roll_2_16 => fifo_out_roll(2*NCALOFIFOS+16),
                     fifo_out_roll_2_17 => fifo_out_roll(2*NCALOFIFOS+17),
                     fifo_out_roll_2_18 => fifo_out_roll(2*NCALOFIFOS+18),
                     fifo_out_roll_2_19 => fifo_out_roll(2*NCALOFIFOS+19)
                 );

        merge2_slice : entity work.calo_router_merge2_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     fifo_out_0_0_pt_V  => fifo_out(0*NCALOFIFOS+ 0).pt,
                     fifo_out_0_1_pt_V  => fifo_out(0*NCALOFIFOS+ 1).pt,
                     fifo_out_0_2_pt_V  => fifo_out(0*NCALOFIFOS+ 2).pt,
                     fifo_out_0_3_pt_V  => fifo_out(0*NCALOFIFOS+ 3).pt,
                     fifo_out_0_4_pt_V  => fifo_out(0*NCALOFIFOS+ 4).pt,
                     fifo_out_0_5_pt_V  => fifo_out(0*NCALOFIFOS+ 5).pt,
                     fifo_out_0_6_pt_V  => fifo_out(0*NCALOFIFOS+ 6).pt,
                     fifo_out_0_7_pt_V  => fifo_out(0*NCALOFIFOS+ 7).pt,
                     fifo_out_0_8_pt_V  => fifo_out(0*NCALOFIFOS+ 8).pt,
                     fifo_out_0_9_pt_V  => fifo_out(0*NCALOFIFOS+ 9).pt,
                     fifo_out_0_10_pt_V => fifo_out(0*NCALOFIFOS+10).pt,
                     fifo_out_0_11_pt_V => fifo_out(0*NCALOFIFOS+11).pt,
                     fifo_out_0_12_pt_V => fifo_out(0*NCALOFIFOS+12).pt,
                     fifo_out_0_13_pt_V => fifo_out(0*NCALOFIFOS+13).pt,
                     fifo_out_0_14_pt_V => fifo_out(0*NCALOFIFOS+14).pt,
                     fifo_out_0_15_pt_V => fifo_out(0*NCALOFIFOS+15).pt,
                     fifo_out_0_16_pt_V => fifo_out(0*NCALOFIFOS+16).pt,
                     fifo_out_0_17_pt_V => fifo_out(0*NCALOFIFOS+17).pt,
                     fifo_out_0_18_pt_V => fifo_out(0*NCALOFIFOS+18).pt,
                     fifo_out_0_19_pt_V => fifo_out(0*NCALOFIFOS+19).pt,
                     fifo_out_1_0_pt_V  => fifo_out(1*NCALOFIFOS+ 0).pt,
                     fifo_out_1_1_pt_V  => fifo_out(1*NCALOFIFOS+ 1).pt,
                     fifo_out_1_2_pt_V  => fifo_out(1*NCALOFIFOS+ 2).pt,
                     fifo_out_1_3_pt_V  => fifo_out(1*NCALOFIFOS+ 3).pt,
                     fifo_out_1_4_pt_V  => fifo_out(1*NCALOFIFOS+ 4).pt,
                     fifo_out_1_5_pt_V  => fifo_out(1*NCALOFIFOS+ 5).pt,
                     fifo_out_1_6_pt_V  => fifo_out(1*NCALOFIFOS+ 6).pt,
                     fifo_out_1_7_pt_V  => fifo_out(1*NCALOFIFOS+ 7).pt,
                     fifo_out_1_8_pt_V  => fifo_out(1*NCALOFIFOS+ 8).pt,
                     fifo_out_1_9_pt_V  => fifo_out(1*NCALOFIFOS+ 9).pt,
                     fifo_out_1_10_pt_V => fifo_out(1*NCALOFIFOS+10).pt,
                     fifo_out_1_11_pt_V => fifo_out(1*NCALOFIFOS+11).pt,
                     fifo_out_1_12_pt_V => fifo_out(1*NCALOFIFOS+12).pt,
                     fifo_out_1_13_pt_V => fifo_out(1*NCALOFIFOS+13).pt,
                     fifo_out_1_14_pt_V => fifo_out(1*NCALOFIFOS+14).pt,
                     fifo_out_1_15_pt_V => fifo_out(1*NCALOFIFOS+15).pt,
                     fifo_out_1_16_pt_V => fifo_out(1*NCALOFIFOS+16).pt,
                     fifo_out_1_17_pt_V => fifo_out(1*NCALOFIFOS+17).pt,
                     fifo_out_1_18_pt_V => fifo_out(1*NCALOFIFOS+18).pt,
                     fifo_out_1_19_pt_V => fifo_out(1*NCALOFIFOS+19).pt,
                     fifo_out_2_0_pt_V  => fifo_out(2*NCALOFIFOS+ 0).pt,
                     fifo_out_2_1_pt_V  => fifo_out(2*NCALOFIFOS+ 1).pt,
                     fifo_out_2_2_pt_V  => fifo_out(2*NCALOFIFOS+ 2).pt,
                     fifo_out_2_3_pt_V  => fifo_out(2*NCALOFIFOS+ 3).pt,
                     fifo_out_2_4_pt_V  => fifo_out(2*NCALOFIFOS+ 4).pt,
                     fifo_out_2_5_pt_V  => fifo_out(2*NCALOFIFOS+ 5).pt,
                     fifo_out_2_6_pt_V  => fifo_out(2*NCALOFIFOS+ 6).pt,
                     fifo_out_2_7_pt_V  => fifo_out(2*NCALOFIFOS+ 7).pt,
                     fifo_out_2_8_pt_V  => fifo_out(2*NCALOFIFOS+ 8).pt,
                     fifo_out_2_9_pt_V  => fifo_out(2*NCALOFIFOS+ 9).pt,
                     fifo_out_2_10_pt_V => fifo_out(2*NCALOFIFOS+10).pt,
                     fifo_out_2_11_pt_V => fifo_out(2*NCALOFIFOS+11).pt,
                     fifo_out_2_12_pt_V => fifo_out(2*NCALOFIFOS+12).pt,
                     fifo_out_2_13_pt_V => fifo_out(2*NCALOFIFOS+13).pt,
                     fifo_out_2_14_pt_V => fifo_out(2*NCALOFIFOS+14).pt,
                     fifo_out_2_15_pt_V => fifo_out(2*NCALOFIFOS+15).pt,
                     fifo_out_2_16_pt_V => fifo_out(2*NCALOFIFOS+16).pt,
                     fifo_out_2_17_pt_V => fifo_out(2*NCALOFIFOS+17).pt,
                     fifo_out_2_18_pt_V => fifo_out(2*NCALOFIFOS+18).pt,
                     fifo_out_2_19_pt_V => fifo_out(2*NCALOFIFOS+19).pt,
                     fifo_out_0_0_eta_V  => fifo_out(0*NCALOFIFOS+ 0).eta,
                     fifo_out_0_1_eta_V  => fifo_out(0*NCALOFIFOS+ 1).eta,
                     fifo_out_0_2_eta_V  => fifo_out(0*NCALOFIFOS+ 2).eta,
                     fifo_out_0_3_eta_V  => fifo_out(0*NCALOFIFOS+ 3).eta,
                     fifo_out_0_4_eta_V  => fifo_out(0*NCALOFIFOS+ 4).eta,
                     fifo_out_0_5_eta_V  => fifo_out(0*NCALOFIFOS+ 5).eta,
                     fifo_out_0_6_eta_V  => fifo_out(0*NCALOFIFOS+ 6).eta,
                     fifo_out_0_7_eta_V  => fifo_out(0*NCALOFIFOS+ 7).eta,
                     fifo_out_0_8_eta_V  => fifo_out(0*NCALOFIFOS+ 8).eta,
                     fifo_out_0_9_eta_V  => fifo_out(0*NCALOFIFOS+ 9).eta,
                     fifo_out_0_10_eta_V => fifo_out(0*NCALOFIFOS+10).eta,
                     fifo_out_0_11_eta_V => fifo_out(0*NCALOFIFOS+11).eta,
                     fifo_out_0_12_eta_V => fifo_out(0*NCALOFIFOS+12).eta,
                     fifo_out_0_13_eta_V => fifo_out(0*NCALOFIFOS+13).eta,
                     fifo_out_0_14_eta_V => fifo_out(0*NCALOFIFOS+14).eta,
                     fifo_out_0_15_eta_V => fifo_out(0*NCALOFIFOS+15).eta,
                     fifo_out_0_16_eta_V => fifo_out(0*NCALOFIFOS+16).eta,
                     fifo_out_0_17_eta_V => fifo_out(0*NCALOFIFOS+17).eta,
                     fifo_out_0_18_eta_V => fifo_out(0*NCALOFIFOS+18).eta,
                     fifo_out_0_19_eta_V => fifo_out(0*NCALOFIFOS+19).eta,
                     fifo_out_1_0_eta_V  => fifo_out(1*NCALOFIFOS+ 0).eta,
                     fifo_out_1_1_eta_V  => fifo_out(1*NCALOFIFOS+ 1).eta,
                     fifo_out_1_2_eta_V  => fifo_out(1*NCALOFIFOS+ 2).eta,
                     fifo_out_1_3_eta_V  => fifo_out(1*NCALOFIFOS+ 3).eta,
                     fifo_out_1_4_eta_V  => fifo_out(1*NCALOFIFOS+ 4).eta,
                     fifo_out_1_5_eta_V  => fifo_out(1*NCALOFIFOS+ 5).eta,
                     fifo_out_1_6_eta_V  => fifo_out(1*NCALOFIFOS+ 6).eta,
                     fifo_out_1_7_eta_V  => fifo_out(1*NCALOFIFOS+ 7).eta,
                     fifo_out_1_8_eta_V  => fifo_out(1*NCALOFIFOS+ 8).eta,
                     fifo_out_1_9_eta_V  => fifo_out(1*NCALOFIFOS+ 9).eta,
                     fifo_out_1_10_eta_V => fifo_out(1*NCALOFIFOS+10).eta,
                     fifo_out_1_11_eta_V => fifo_out(1*NCALOFIFOS+11).eta,
                     fifo_out_1_12_eta_V => fifo_out(1*NCALOFIFOS+12).eta,
                     fifo_out_1_13_eta_V => fifo_out(1*NCALOFIFOS+13).eta,
                     fifo_out_1_14_eta_V => fifo_out(1*NCALOFIFOS+14).eta,
                     fifo_out_1_15_eta_V => fifo_out(1*NCALOFIFOS+15).eta,
                     fifo_out_1_16_eta_V => fifo_out(1*NCALOFIFOS+16).eta,
                     fifo_out_1_17_eta_V => fifo_out(1*NCALOFIFOS+17).eta,
                     fifo_out_1_18_eta_V => fifo_out(1*NCALOFIFOS+18).eta,
                     fifo_out_1_19_eta_V => fifo_out(1*NCALOFIFOS+19).eta,
                     fifo_out_2_0_eta_V  => fifo_out(2*NCALOFIFOS+ 0).eta,
                     fifo_out_2_1_eta_V  => fifo_out(2*NCALOFIFOS+ 1).eta,
                     fifo_out_2_2_eta_V  => fifo_out(2*NCALOFIFOS+ 2).eta,
                     fifo_out_2_3_eta_V  => fifo_out(2*NCALOFIFOS+ 3).eta,
                     fifo_out_2_4_eta_V  => fifo_out(2*NCALOFIFOS+ 4).eta,
                     fifo_out_2_5_eta_V  => fifo_out(2*NCALOFIFOS+ 5).eta,
                     fifo_out_2_6_eta_V  => fifo_out(2*NCALOFIFOS+ 6).eta,
                     fifo_out_2_7_eta_V  => fifo_out(2*NCALOFIFOS+ 7).eta,
                     fifo_out_2_8_eta_V  => fifo_out(2*NCALOFIFOS+ 8).eta,
                     fifo_out_2_9_eta_V  => fifo_out(2*NCALOFIFOS+ 9).eta,
                     fifo_out_2_10_eta_V => fifo_out(2*NCALOFIFOS+10).eta,
                     fifo_out_2_11_eta_V => fifo_out(2*NCALOFIFOS+11).eta,
                     fifo_out_2_12_eta_V => fifo_out(2*NCALOFIFOS+12).eta,
                     fifo_out_2_13_eta_V => fifo_out(2*NCALOFIFOS+13).eta,
                     fifo_out_2_14_eta_V => fifo_out(2*NCALOFIFOS+14).eta,
                     fifo_out_2_15_eta_V => fifo_out(2*NCALOFIFOS+15).eta,
                     fifo_out_2_16_eta_V => fifo_out(2*NCALOFIFOS+16).eta,
                     fifo_out_2_17_eta_V => fifo_out(2*NCALOFIFOS+17).eta,
                     fifo_out_2_18_eta_V => fifo_out(2*NCALOFIFOS+18).eta,
                     fifo_out_2_19_eta_V => fifo_out(2*NCALOFIFOS+19).eta,
                     fifo_out_0_0_phi_V  => fifo_out(0*NCALOFIFOS+ 0).phi,
                     fifo_out_0_1_phi_V  => fifo_out(0*NCALOFIFOS+ 1).phi,
                     fifo_out_0_2_phi_V  => fifo_out(0*NCALOFIFOS+ 2).phi,
                     fifo_out_0_3_phi_V  => fifo_out(0*NCALOFIFOS+ 3).phi,
                     fifo_out_0_4_phi_V  => fifo_out(0*NCALOFIFOS+ 4).phi,
                     fifo_out_0_5_phi_V  => fifo_out(0*NCALOFIFOS+ 5).phi,
                     fifo_out_0_6_phi_V  => fifo_out(0*NCALOFIFOS+ 6).phi,
                     fifo_out_0_7_phi_V  => fifo_out(0*NCALOFIFOS+ 7).phi,
                     fifo_out_0_8_phi_V  => fifo_out(0*NCALOFIFOS+ 8).phi,
                     fifo_out_0_9_phi_V  => fifo_out(0*NCALOFIFOS+ 9).phi,
                     fifo_out_0_10_phi_V => fifo_out(0*NCALOFIFOS+10).phi,
                     fifo_out_0_11_phi_V => fifo_out(0*NCALOFIFOS+11).phi,
                     fifo_out_0_12_phi_V => fifo_out(0*NCALOFIFOS+12).phi,
                     fifo_out_0_13_phi_V => fifo_out(0*NCALOFIFOS+13).phi,
                     fifo_out_0_14_phi_V => fifo_out(0*NCALOFIFOS+14).phi,
                     fifo_out_0_15_phi_V => fifo_out(0*NCALOFIFOS+15).phi,
                     fifo_out_0_16_phi_V => fifo_out(0*NCALOFIFOS+16).phi,
                     fifo_out_0_17_phi_V => fifo_out(0*NCALOFIFOS+17).phi,
                     fifo_out_0_18_phi_V => fifo_out(0*NCALOFIFOS+18).phi,
                     fifo_out_0_19_phi_V => fifo_out(0*NCALOFIFOS+19).phi,
                     fifo_out_1_0_phi_V  => fifo_out(1*NCALOFIFOS+ 0).phi,
                     fifo_out_1_1_phi_V  => fifo_out(1*NCALOFIFOS+ 1).phi,
                     fifo_out_1_2_phi_V  => fifo_out(1*NCALOFIFOS+ 2).phi,
                     fifo_out_1_3_phi_V  => fifo_out(1*NCALOFIFOS+ 3).phi,
                     fifo_out_1_4_phi_V  => fifo_out(1*NCALOFIFOS+ 4).phi,
                     fifo_out_1_5_phi_V  => fifo_out(1*NCALOFIFOS+ 5).phi,
                     fifo_out_1_6_phi_V  => fifo_out(1*NCALOFIFOS+ 6).phi,
                     fifo_out_1_7_phi_V  => fifo_out(1*NCALOFIFOS+ 7).phi,
                     fifo_out_1_8_phi_V  => fifo_out(1*NCALOFIFOS+ 8).phi,
                     fifo_out_1_9_phi_V  => fifo_out(1*NCALOFIFOS+ 9).phi,
                     fifo_out_1_10_phi_V => fifo_out(1*NCALOFIFOS+10).phi,
                     fifo_out_1_11_phi_V => fifo_out(1*NCALOFIFOS+11).phi,
                     fifo_out_1_12_phi_V => fifo_out(1*NCALOFIFOS+12).phi,
                     fifo_out_1_13_phi_V => fifo_out(1*NCALOFIFOS+13).phi,
                     fifo_out_1_14_phi_V => fifo_out(1*NCALOFIFOS+14).phi,
                     fifo_out_1_15_phi_V => fifo_out(1*NCALOFIFOS+15).phi,
                     fifo_out_1_16_phi_V => fifo_out(1*NCALOFIFOS+16).phi,
                     fifo_out_1_17_phi_V => fifo_out(1*NCALOFIFOS+17).phi,
                     fifo_out_1_18_phi_V => fifo_out(1*NCALOFIFOS+18).phi,
                     fifo_out_1_19_phi_V => fifo_out(1*NCALOFIFOS+19).phi,
                     fifo_out_2_0_phi_V  => fifo_out(2*NCALOFIFOS+ 0).phi,
                     fifo_out_2_1_phi_V  => fifo_out(2*NCALOFIFOS+ 1).phi,
                     fifo_out_2_2_phi_V  => fifo_out(2*NCALOFIFOS+ 2).phi,
                     fifo_out_2_3_phi_V  => fifo_out(2*NCALOFIFOS+ 3).phi,
                     fifo_out_2_4_phi_V  => fifo_out(2*NCALOFIFOS+ 4).phi,
                     fifo_out_2_5_phi_V  => fifo_out(2*NCALOFIFOS+ 5).phi,
                     fifo_out_2_6_phi_V  => fifo_out(2*NCALOFIFOS+ 6).phi,
                     fifo_out_2_7_phi_V  => fifo_out(2*NCALOFIFOS+ 7).phi,
                     fifo_out_2_8_phi_V  => fifo_out(2*NCALOFIFOS+ 8).phi,
                     fifo_out_2_9_phi_V  => fifo_out(2*NCALOFIFOS+ 9).phi,
                     fifo_out_2_10_phi_V => fifo_out(2*NCALOFIFOS+10).phi,
                     fifo_out_2_11_phi_V => fifo_out(2*NCALOFIFOS+11).phi,
                     fifo_out_2_12_phi_V => fifo_out(2*NCALOFIFOS+12).phi,
                     fifo_out_2_13_phi_V => fifo_out(2*NCALOFIFOS+13).phi,
                     fifo_out_2_14_phi_V => fifo_out(2*NCALOFIFOS+14).phi,
                     fifo_out_2_15_phi_V => fifo_out(2*NCALOFIFOS+15).phi,
                     fifo_out_2_16_phi_V => fifo_out(2*NCALOFIFOS+16).phi,
                     fifo_out_2_17_phi_V => fifo_out(2*NCALOFIFOS+17).phi,
                     fifo_out_2_18_phi_V => fifo_out(2*NCALOFIFOS+18).phi,
                     fifo_out_2_19_phi_V => fifo_out(2*NCALOFIFOS+19).phi,
                     fifo_out_0_0_rest_V  => fifo_out(0*NCALOFIFOS+ 0).rest,
                     fifo_out_0_1_rest_V  => fifo_out(0*NCALOFIFOS+ 1).rest,
                     fifo_out_0_2_rest_V  => fifo_out(0*NCALOFIFOS+ 2).rest,
                     fifo_out_0_3_rest_V  => fifo_out(0*NCALOFIFOS+ 3).rest,
                     fifo_out_0_4_rest_V  => fifo_out(0*NCALOFIFOS+ 4).rest,
                     fifo_out_0_5_rest_V  => fifo_out(0*NCALOFIFOS+ 5).rest,
                     fifo_out_0_6_rest_V  => fifo_out(0*NCALOFIFOS+ 6).rest,
                     fifo_out_0_7_rest_V  => fifo_out(0*NCALOFIFOS+ 7).rest,
                     fifo_out_0_8_rest_V  => fifo_out(0*NCALOFIFOS+ 8).rest,
                     fifo_out_0_9_rest_V  => fifo_out(0*NCALOFIFOS+ 9).rest,
                     fifo_out_0_10_rest_V => fifo_out(0*NCALOFIFOS+10).rest,
                     fifo_out_0_11_rest_V => fifo_out(0*NCALOFIFOS+11).rest,
                     fifo_out_0_12_rest_V => fifo_out(0*NCALOFIFOS+12).rest,
                     fifo_out_0_13_rest_V => fifo_out(0*NCALOFIFOS+13).rest,
                     fifo_out_0_14_rest_V => fifo_out(0*NCALOFIFOS+14).rest,
                     fifo_out_0_15_rest_V => fifo_out(0*NCALOFIFOS+15).rest,
                     fifo_out_0_16_rest_V => fifo_out(0*NCALOFIFOS+16).rest,
                     fifo_out_0_17_rest_V => fifo_out(0*NCALOFIFOS+17).rest,
                     fifo_out_0_18_rest_V => fifo_out(0*NCALOFIFOS+18).rest,
                     fifo_out_0_19_rest_V => fifo_out(0*NCALOFIFOS+19).rest,
                     fifo_out_1_0_rest_V  => fifo_out(1*NCALOFIFOS+ 0).rest,
                     fifo_out_1_1_rest_V  => fifo_out(1*NCALOFIFOS+ 1).rest,
                     fifo_out_1_2_rest_V  => fifo_out(1*NCALOFIFOS+ 2).rest,
                     fifo_out_1_3_rest_V  => fifo_out(1*NCALOFIFOS+ 3).rest,
                     fifo_out_1_4_rest_V  => fifo_out(1*NCALOFIFOS+ 4).rest,
                     fifo_out_1_5_rest_V  => fifo_out(1*NCALOFIFOS+ 5).rest,
                     fifo_out_1_6_rest_V  => fifo_out(1*NCALOFIFOS+ 6).rest,
                     fifo_out_1_7_rest_V  => fifo_out(1*NCALOFIFOS+ 7).rest,
                     fifo_out_1_8_rest_V  => fifo_out(1*NCALOFIFOS+ 8).rest,
                     fifo_out_1_9_rest_V  => fifo_out(1*NCALOFIFOS+ 9).rest,
                     fifo_out_1_10_rest_V => fifo_out(1*NCALOFIFOS+10).rest,
                     fifo_out_1_11_rest_V => fifo_out(1*NCALOFIFOS+11).rest,
                     fifo_out_1_12_rest_V => fifo_out(1*NCALOFIFOS+12).rest,
                     fifo_out_1_13_rest_V => fifo_out(1*NCALOFIFOS+13).rest,
                     fifo_out_1_14_rest_V => fifo_out(1*NCALOFIFOS+14).rest,
                     fifo_out_1_15_rest_V => fifo_out(1*NCALOFIFOS+15).rest,
                     fifo_out_1_16_rest_V => fifo_out(1*NCALOFIFOS+16).rest,
                     fifo_out_1_17_rest_V => fifo_out(1*NCALOFIFOS+17).rest,
                     fifo_out_1_18_rest_V => fifo_out(1*NCALOFIFOS+18).rest,
                     fifo_out_1_19_rest_V => fifo_out(1*NCALOFIFOS+19).rest,
                     fifo_out_2_0_rest_V  => fifo_out(2*NCALOFIFOS+ 0).rest,
                     fifo_out_2_1_rest_V  => fifo_out(2*NCALOFIFOS+ 1).rest,
                     fifo_out_2_2_rest_V  => fifo_out(2*NCALOFIFOS+ 2).rest,
                     fifo_out_2_3_rest_V  => fifo_out(2*NCALOFIFOS+ 3).rest,
                     fifo_out_2_4_rest_V  => fifo_out(2*NCALOFIFOS+ 4).rest,
                     fifo_out_2_5_rest_V  => fifo_out(2*NCALOFIFOS+ 5).rest,
                     fifo_out_2_6_rest_V  => fifo_out(2*NCALOFIFOS+ 6).rest,
                     fifo_out_2_7_rest_V  => fifo_out(2*NCALOFIFOS+ 7).rest,
                     fifo_out_2_8_rest_V  => fifo_out(2*NCALOFIFOS+ 8).rest,
                     fifo_out_2_9_rest_V  => fifo_out(2*NCALOFIFOS+ 9).rest,
                     fifo_out_2_10_rest_V => fifo_out(2*NCALOFIFOS+10).rest,
                     fifo_out_2_11_rest_V => fifo_out(2*NCALOFIFOS+11).rest,
                     fifo_out_2_12_rest_V => fifo_out(2*NCALOFIFOS+12).rest,
                     fifo_out_2_13_rest_V => fifo_out(2*NCALOFIFOS+13).rest,
                     fifo_out_2_14_rest_V => fifo_out(2*NCALOFIFOS+14).rest,
                     fifo_out_2_15_rest_V => fifo_out(2*NCALOFIFOS+15).rest,
                     fifo_out_2_16_rest_V => fifo_out(2*NCALOFIFOS+16).rest,
                     fifo_out_2_17_rest_V => fifo_out(2*NCALOFIFOS+17).rest,
                     fifo_out_2_18_rest_V => fifo_out(2*NCALOFIFOS+18).rest,
                     fifo_out_2_19_rest_V => fifo_out(2*NCALOFIFOS+19).rest,
                     fifo_full_0_0  => fifo_full(0*NCALOFIFOS+ 0),
                     fifo_full_0_1  => fifo_full(0*NCALOFIFOS+ 1),
                     fifo_full_0_2  => fifo_full(0*NCALOFIFOS+ 2),
                     fifo_full_0_3  => fifo_full(0*NCALOFIFOS+ 3),
                     fifo_full_0_4  => fifo_full(0*NCALOFIFOS+ 4),
                     fifo_full_0_5  => fifo_full(0*NCALOFIFOS+ 5),
                     fifo_full_0_6  => fifo_full(0*NCALOFIFOS+ 6),
                     fifo_full_0_7  => fifo_full(0*NCALOFIFOS+ 7),
                     fifo_full_0_8  => fifo_full(0*NCALOFIFOS+ 8),
                     fifo_full_0_9  => fifo_full(0*NCALOFIFOS+ 9),
                     fifo_full_0_10 => fifo_full(0*NCALOFIFOS+10),
                     fifo_full_0_11 => fifo_full(0*NCALOFIFOS+11),
                     fifo_full_0_12 => fifo_full(0*NCALOFIFOS+12),
                     fifo_full_0_13 => fifo_full(0*NCALOFIFOS+13),
                     fifo_full_0_14 => fifo_full(0*NCALOFIFOS+14),
                     fifo_full_0_15 => fifo_full(0*NCALOFIFOS+15),
                     fifo_full_0_16 => fifo_full(0*NCALOFIFOS+16),
                     fifo_full_0_17 => fifo_full(0*NCALOFIFOS+17),
                     fifo_full_0_18 => fifo_full(0*NCALOFIFOS+18),
                     fifo_full_0_19 => fifo_full(0*NCALOFIFOS+19),
                     fifo_full_1_0  => fifo_full(1*NCALOFIFOS+ 0),
                     fifo_full_1_1  => fifo_full(1*NCALOFIFOS+ 1),
                     fifo_full_1_2  => fifo_full(1*NCALOFIFOS+ 2),
                     fifo_full_1_3  => fifo_full(1*NCALOFIFOS+ 3),
                     fifo_full_1_4  => fifo_full(1*NCALOFIFOS+ 4),
                     fifo_full_1_5  => fifo_full(1*NCALOFIFOS+ 5),
                     fifo_full_1_6  => fifo_full(1*NCALOFIFOS+ 6),
                     fifo_full_1_7  => fifo_full(1*NCALOFIFOS+ 7),
                     fifo_full_1_8  => fifo_full(1*NCALOFIFOS+ 8),
                     fifo_full_1_9  => fifo_full(1*NCALOFIFOS+ 9),
                     fifo_full_1_10 => fifo_full(1*NCALOFIFOS+10),
                     fifo_full_1_11 => fifo_full(1*NCALOFIFOS+11),
                     fifo_full_1_12 => fifo_full(1*NCALOFIFOS+12),
                     fifo_full_1_13 => fifo_full(1*NCALOFIFOS+13),
                     fifo_full_1_14 => fifo_full(1*NCALOFIFOS+14),
                     fifo_full_1_15 => fifo_full(1*NCALOFIFOS+15),
                     fifo_full_1_16 => fifo_full(1*NCALOFIFOS+16),
                     fifo_full_1_17 => fifo_full(1*NCALOFIFOS+17),
                     fifo_full_1_18 => fifo_full(1*NCALOFIFOS+18),
                     fifo_full_1_19 => fifo_full(1*NCALOFIFOS+19),
                     fifo_full_2_0  => fifo_full(2*NCALOFIFOS+ 0),
                     fifo_full_2_1  => fifo_full(2*NCALOFIFOS+ 1),
                     fifo_full_2_2  => fifo_full(2*NCALOFIFOS+ 2),
                     fifo_full_2_3  => fifo_full(2*NCALOFIFOS+ 3),
                     fifo_full_2_4  => fifo_full(2*NCALOFIFOS+ 4),
                     fifo_full_2_5  => fifo_full(2*NCALOFIFOS+ 5),
                     fifo_full_2_6  => fifo_full(2*NCALOFIFOS+ 6),
                     fifo_full_2_7  => fifo_full(2*NCALOFIFOS+ 7),
                     fifo_full_2_8  => fifo_full(2*NCALOFIFOS+ 8),
                     fifo_full_2_9  => fifo_full(2*NCALOFIFOS+ 9),
                     fifo_full_2_10 => fifo_full(2*NCALOFIFOS+10),
                     fifo_full_2_11 => fifo_full(2*NCALOFIFOS+11),
                     fifo_full_2_12 => fifo_full(2*NCALOFIFOS+12),
                     fifo_full_2_13 => fifo_full(2*NCALOFIFOS+13),
                     fifo_full_2_14 => fifo_full(2*NCALOFIFOS+14),
                     fifo_full_2_15 => fifo_full(2*NCALOFIFOS+15),
                     fifo_full_2_16 => fifo_full(2*NCALOFIFOS+16),
                     fifo_full_2_17 => fifo_full(2*NCALOFIFOS+17),
                     fifo_full_2_18 => fifo_full(2*NCALOFIFOS+18),
                     fifo_full_2_19 => fifo_full(2*NCALOFIFOS+19),
                     fifo_out_valid_0_0  => fifo_out_valid(0*NCALOFIFOS+ 0),
                     fifo_out_valid_0_1  => fifo_out_valid(0*NCALOFIFOS+ 1),
                     fifo_out_valid_0_2  => fifo_out_valid(0*NCALOFIFOS+ 2),
                     fifo_out_valid_0_3  => fifo_out_valid(0*NCALOFIFOS+ 3),
                     fifo_out_valid_0_4  => fifo_out_valid(0*NCALOFIFOS+ 4),
                     fifo_out_valid_0_5  => fifo_out_valid(0*NCALOFIFOS+ 5),
                     fifo_out_valid_0_6  => fifo_out_valid(0*NCALOFIFOS+ 6),
                     fifo_out_valid_0_7  => fifo_out_valid(0*NCALOFIFOS+ 7),
                     fifo_out_valid_0_8  => fifo_out_valid(0*NCALOFIFOS+ 8),
                     fifo_out_valid_0_9  => fifo_out_valid(0*NCALOFIFOS+ 9),
                     fifo_out_valid_0_10 => fifo_out_valid(0*NCALOFIFOS+10),
                     fifo_out_valid_0_11 => fifo_out_valid(0*NCALOFIFOS+11),
                     fifo_out_valid_0_12 => fifo_out_valid(0*NCALOFIFOS+12),
                     fifo_out_valid_0_13 => fifo_out_valid(0*NCALOFIFOS+13),
                     fifo_out_valid_0_14 => fifo_out_valid(0*NCALOFIFOS+14),
                     fifo_out_valid_0_15 => fifo_out_valid(0*NCALOFIFOS+15),
                     fifo_out_valid_0_16 => fifo_out_valid(0*NCALOFIFOS+16),
                     fifo_out_valid_0_17 => fifo_out_valid(0*NCALOFIFOS+17),
                     fifo_out_valid_0_18 => fifo_out_valid(0*NCALOFIFOS+18),
                     fifo_out_valid_0_19 => fifo_out_valid(0*NCALOFIFOS+19),
                     fifo_out_valid_1_0  => fifo_out_valid(1*NCALOFIFOS+ 0),
                     fifo_out_valid_1_1  => fifo_out_valid(1*NCALOFIFOS+ 1),
                     fifo_out_valid_1_2  => fifo_out_valid(1*NCALOFIFOS+ 2),
                     fifo_out_valid_1_3  => fifo_out_valid(1*NCALOFIFOS+ 3),
                     fifo_out_valid_1_4  => fifo_out_valid(1*NCALOFIFOS+ 4),
                     fifo_out_valid_1_5  => fifo_out_valid(1*NCALOFIFOS+ 5),
                     fifo_out_valid_1_6  => fifo_out_valid(1*NCALOFIFOS+ 6),
                     fifo_out_valid_1_7  => fifo_out_valid(1*NCALOFIFOS+ 7),
                     fifo_out_valid_1_8  => fifo_out_valid(1*NCALOFIFOS+ 8),
                     fifo_out_valid_1_9  => fifo_out_valid(1*NCALOFIFOS+ 9),
                     fifo_out_valid_1_10 => fifo_out_valid(1*NCALOFIFOS+10),
                     fifo_out_valid_1_11 => fifo_out_valid(1*NCALOFIFOS+11),
                     fifo_out_valid_1_12 => fifo_out_valid(1*NCALOFIFOS+12),
                     fifo_out_valid_1_13 => fifo_out_valid(1*NCALOFIFOS+13),
                     fifo_out_valid_1_14 => fifo_out_valid(1*NCALOFIFOS+14),
                     fifo_out_valid_1_15 => fifo_out_valid(1*NCALOFIFOS+15),
                     fifo_out_valid_1_16 => fifo_out_valid(1*NCALOFIFOS+16),
                     fifo_out_valid_1_17 => fifo_out_valid(1*NCALOFIFOS+17),
                     fifo_out_valid_1_18 => fifo_out_valid(1*NCALOFIFOS+18),
                     fifo_out_valid_1_19 => fifo_out_valid(1*NCALOFIFOS+19),
                     fifo_out_valid_2_0  => fifo_out_valid(2*NCALOFIFOS+ 0),
                     fifo_out_valid_2_1  => fifo_out_valid(2*NCALOFIFOS+ 1),
                     fifo_out_valid_2_2  => fifo_out_valid(2*NCALOFIFOS+ 2),
                     fifo_out_valid_2_3  => fifo_out_valid(2*NCALOFIFOS+ 3),
                     fifo_out_valid_2_4  => fifo_out_valid(2*NCALOFIFOS+ 4),
                     fifo_out_valid_2_5  => fifo_out_valid(2*NCALOFIFOS+ 5),
                     fifo_out_valid_2_6  => fifo_out_valid(2*NCALOFIFOS+ 6),
                     fifo_out_valid_2_7  => fifo_out_valid(2*NCALOFIFOS+ 7),
                     fifo_out_valid_2_8  => fifo_out_valid(2*NCALOFIFOS+ 8),
                     fifo_out_valid_2_9  => fifo_out_valid(2*NCALOFIFOS+ 9),
                     fifo_out_valid_2_10 => fifo_out_valid(2*NCALOFIFOS+10),
                     fifo_out_valid_2_11 => fifo_out_valid(2*NCALOFIFOS+11),
                     fifo_out_valid_2_12 => fifo_out_valid(2*NCALOFIFOS+12),
                     fifo_out_valid_2_13 => fifo_out_valid(2*NCALOFIFOS+13),
                     fifo_out_valid_2_14 => fifo_out_valid(2*NCALOFIFOS+14),
                     fifo_out_valid_2_15 => fifo_out_valid(2*NCALOFIFOS+15),
                     fifo_out_valid_2_16 => fifo_out_valid(2*NCALOFIFOS+16),
                     fifo_out_valid_2_17 => fifo_out_valid(2*NCALOFIFOS+17),
                     fifo_out_valid_2_18 => fifo_out_valid(2*NCALOFIFOS+18),
                     fifo_out_valid_2_19 => fifo_out_valid(2*NCALOFIFOS+19),
                     fifo_out_roll_0_0  => fifo_out_roll(0*NCALOFIFOS+ 0),
                     fifo_out_roll_0_1  => fifo_out_roll(0*NCALOFIFOS+ 1),
                     fifo_out_roll_0_2  => fifo_out_roll(0*NCALOFIFOS+ 2),
                     fifo_out_roll_0_3  => fifo_out_roll(0*NCALOFIFOS+ 3),
                     fifo_out_roll_0_4  => fifo_out_roll(0*NCALOFIFOS+ 4),
                     fifo_out_roll_0_5  => fifo_out_roll(0*NCALOFIFOS+ 5),
                     fifo_out_roll_0_6  => fifo_out_roll(0*NCALOFIFOS+ 6),
                     fifo_out_roll_0_7  => fifo_out_roll(0*NCALOFIFOS+ 7),
                     fifo_out_roll_0_8  => fifo_out_roll(0*NCALOFIFOS+ 8),
                     fifo_out_roll_0_9  => fifo_out_roll(0*NCALOFIFOS+ 9),
                     fifo_out_roll_0_10 => fifo_out_roll(0*NCALOFIFOS+10),
                     fifo_out_roll_0_11 => fifo_out_roll(0*NCALOFIFOS+11),
                     fifo_out_roll_0_12 => fifo_out_roll(0*NCALOFIFOS+12),
                     fifo_out_roll_0_13 => fifo_out_roll(0*NCALOFIFOS+13),
                     fifo_out_roll_0_14 => fifo_out_roll(0*NCALOFIFOS+14),
                     fifo_out_roll_0_15 => fifo_out_roll(0*NCALOFIFOS+15),
                     fifo_out_roll_0_16 => fifo_out_roll(0*NCALOFIFOS+16),
                     fifo_out_roll_0_17 => fifo_out_roll(0*NCALOFIFOS+17),
                     fifo_out_roll_0_18 => fifo_out_roll(0*NCALOFIFOS+18),
                     fifo_out_roll_0_19 => fifo_out_roll(0*NCALOFIFOS+19),
                     fifo_out_roll_1_0  => fifo_out_roll(1*NCALOFIFOS+ 0),
                     fifo_out_roll_1_1  => fifo_out_roll(1*NCALOFIFOS+ 1),
                     fifo_out_roll_1_2  => fifo_out_roll(1*NCALOFIFOS+ 2),
                     fifo_out_roll_1_3  => fifo_out_roll(1*NCALOFIFOS+ 3),
                     fifo_out_roll_1_4  => fifo_out_roll(1*NCALOFIFOS+ 4),
                     fifo_out_roll_1_5  => fifo_out_roll(1*NCALOFIFOS+ 5),
                     fifo_out_roll_1_6  => fifo_out_roll(1*NCALOFIFOS+ 6),
                     fifo_out_roll_1_7  => fifo_out_roll(1*NCALOFIFOS+ 7),
                     fifo_out_roll_1_8  => fifo_out_roll(1*NCALOFIFOS+ 8),
                     fifo_out_roll_1_9  => fifo_out_roll(1*NCALOFIFOS+ 9),
                     fifo_out_roll_1_10 => fifo_out_roll(1*NCALOFIFOS+10),
                     fifo_out_roll_1_11 => fifo_out_roll(1*NCALOFIFOS+11),
                     fifo_out_roll_1_12 => fifo_out_roll(1*NCALOFIFOS+12),
                     fifo_out_roll_1_13 => fifo_out_roll(1*NCALOFIFOS+13),
                     fifo_out_roll_1_14 => fifo_out_roll(1*NCALOFIFOS+14),
                     fifo_out_roll_1_15 => fifo_out_roll(1*NCALOFIFOS+15),
                     fifo_out_roll_1_16 => fifo_out_roll(1*NCALOFIFOS+16),
                     fifo_out_roll_1_17 => fifo_out_roll(1*NCALOFIFOS+17),
                     fifo_out_roll_1_18 => fifo_out_roll(1*NCALOFIFOS+18),
                     fifo_out_roll_1_19 => fifo_out_roll(1*NCALOFIFOS+19),
                     fifo_out_roll_2_0  => fifo_out_roll(2*NCALOFIFOS+ 0),
                     fifo_out_roll_2_1  => fifo_out_roll(2*NCALOFIFOS+ 1),
                     fifo_out_roll_2_2  => fifo_out_roll(2*NCALOFIFOS+ 2),
                     fifo_out_roll_2_3  => fifo_out_roll(2*NCALOFIFOS+ 3),
                     fifo_out_roll_2_4  => fifo_out_roll(2*NCALOFIFOS+ 4),
                     fifo_out_roll_2_5  => fifo_out_roll(2*NCALOFIFOS+ 5),
                     fifo_out_roll_2_6  => fifo_out_roll(2*NCALOFIFOS+ 6),
                     fifo_out_roll_2_7  => fifo_out_roll(2*NCALOFIFOS+ 7),
                     fifo_out_roll_2_8  => fifo_out_roll(2*NCALOFIFOS+ 8),
                     fifo_out_roll_2_9  => fifo_out_roll(2*NCALOFIFOS+ 9),
                     fifo_out_roll_2_10 => fifo_out_roll(2*NCALOFIFOS+10),
                     fifo_out_roll_2_11 => fifo_out_roll(2*NCALOFIFOS+11),
                     fifo_out_roll_2_12 => fifo_out_roll(2*NCALOFIFOS+12),
                     fifo_out_roll_2_13 => fifo_out_roll(2*NCALOFIFOS+13),
                     fifo_out_roll_2_14 => fifo_out_roll(2*NCALOFIFOS+14),
                     fifo_out_roll_2_15 => fifo_out_roll(2*NCALOFIFOS+15),
                     fifo_out_roll_2_16 => fifo_out_roll(2*NCALOFIFOS+16),
                     fifo_out_roll_2_17 => fifo_out_roll(2*NCALOFIFOS+17),
                     fifo_out_roll_2_18 => fifo_out_roll(2*NCALOFIFOS+18),
                     fifo_out_roll_2_19 => fifo_out_roll(2*NCALOFIFOS+19),
                     merged_out_0_0_pt_V  => merged2_out(0*NCALOFIFOS/2+0).pt,
                     merged_out_0_1_pt_V  => merged2_out(0*NCALOFIFOS/2+1).pt,
                     merged_out_0_2_pt_V  => merged2_out(0*NCALOFIFOS/2+2).pt,
                     merged_out_0_3_pt_V  => merged2_out(0*NCALOFIFOS/2+3).pt,
                     merged_out_0_4_pt_V  => merged2_out(0*NCALOFIFOS/2+4).pt,
                     merged_out_0_5_pt_V  => merged2_out(0*NCALOFIFOS/2+5).pt,
                     merged_out_0_6_pt_V  => merged2_out(0*NCALOFIFOS/2+6).pt,
                     merged_out_0_7_pt_V  => merged2_out(0*NCALOFIFOS/2+7).pt,
                     merged_out_0_8_pt_V  => merged2_out(0*NCALOFIFOS/2+8).pt,
                     merged_out_0_9_pt_V  => merged2_out(0*NCALOFIFOS/2+9).pt,
                     merged_out_1_0_pt_V  => merged2_out(1*NCALOFIFOS/2+0).pt,
                     merged_out_1_1_pt_V  => merged2_out(1*NCALOFIFOS/2+1).pt,
                     merged_out_1_2_pt_V  => merged2_out(1*NCALOFIFOS/2+2).pt,
                     merged_out_1_3_pt_V  => merged2_out(1*NCALOFIFOS/2+3).pt,
                     merged_out_1_4_pt_V  => merged2_out(1*NCALOFIFOS/2+4).pt,
                     merged_out_1_5_pt_V  => merged2_out(1*NCALOFIFOS/2+5).pt,
                     merged_out_1_6_pt_V  => merged2_out(1*NCALOFIFOS/2+6).pt,
                     merged_out_1_7_pt_V  => merged2_out(1*NCALOFIFOS/2+7).pt,
                     merged_out_1_8_pt_V  => merged2_out(1*NCALOFIFOS/2+8).pt,
                     merged_out_1_9_pt_V  => merged2_out(1*NCALOFIFOS/2+9).pt,
                     merged_out_2_0_pt_V  => merged2_out(2*NCALOFIFOS/2+0).pt,
                     merged_out_2_1_pt_V  => merged2_out(2*NCALOFIFOS/2+1).pt,
                     merged_out_2_2_pt_V  => merged2_out(2*NCALOFIFOS/2+2).pt,
                     merged_out_2_3_pt_V  => merged2_out(2*NCALOFIFOS/2+3).pt,
                     merged_out_2_4_pt_V  => merged2_out(2*NCALOFIFOS/2+4).pt,
                     merged_out_2_5_pt_V  => merged2_out(2*NCALOFIFOS/2+5).pt,
                     merged_out_2_6_pt_V  => merged2_out(2*NCALOFIFOS/2+6).pt,
                     merged_out_2_7_pt_V  => merged2_out(2*NCALOFIFOS/2+7).pt,
                     merged_out_2_8_pt_V  => merged2_out(2*NCALOFIFOS/2+8).pt,
                     merged_out_2_9_pt_V  => merged2_out(2*NCALOFIFOS/2+9).pt,
                     merged_out_0_0_eta_V  => merged2_out(0*NCALOFIFOS/2+0).eta,
                     merged_out_0_1_eta_V  => merged2_out(0*NCALOFIFOS/2+1).eta,
                     merged_out_0_2_eta_V  => merged2_out(0*NCALOFIFOS/2+2).eta,
                     merged_out_0_3_eta_V  => merged2_out(0*NCALOFIFOS/2+3).eta,
                     merged_out_0_4_eta_V  => merged2_out(0*NCALOFIFOS/2+4).eta,
                     merged_out_0_5_eta_V  => merged2_out(0*NCALOFIFOS/2+5).eta,
                     merged_out_0_6_eta_V  => merged2_out(0*NCALOFIFOS/2+6).eta,
                     merged_out_0_7_eta_V  => merged2_out(0*NCALOFIFOS/2+7).eta,
                     merged_out_0_8_eta_V  => merged2_out(0*NCALOFIFOS/2+8).eta,
                     merged_out_0_9_eta_V  => merged2_out(0*NCALOFIFOS/2+9).eta,
                     merged_out_1_0_eta_V  => merged2_out(1*NCALOFIFOS/2+0).eta,
                     merged_out_1_1_eta_V  => merged2_out(1*NCALOFIFOS/2+1).eta,
                     merged_out_1_2_eta_V  => merged2_out(1*NCALOFIFOS/2+2).eta,
                     merged_out_1_3_eta_V  => merged2_out(1*NCALOFIFOS/2+3).eta,
                     merged_out_1_4_eta_V  => merged2_out(1*NCALOFIFOS/2+4).eta,
                     merged_out_1_5_eta_V  => merged2_out(1*NCALOFIFOS/2+5).eta,
                     merged_out_1_6_eta_V  => merged2_out(1*NCALOFIFOS/2+6).eta,
                     merged_out_1_7_eta_V  => merged2_out(1*NCALOFIFOS/2+7).eta,
                     merged_out_1_8_eta_V  => merged2_out(1*NCALOFIFOS/2+8).eta,
                     merged_out_1_9_eta_V  => merged2_out(1*NCALOFIFOS/2+9).eta,
                     merged_out_2_0_eta_V  => merged2_out(2*NCALOFIFOS/2+0).eta,
                     merged_out_2_1_eta_V  => merged2_out(2*NCALOFIFOS/2+1).eta,
                     merged_out_2_2_eta_V  => merged2_out(2*NCALOFIFOS/2+2).eta,
                     merged_out_2_3_eta_V  => merged2_out(2*NCALOFIFOS/2+3).eta,
                     merged_out_2_4_eta_V  => merged2_out(2*NCALOFIFOS/2+4).eta,
                     merged_out_2_5_eta_V  => merged2_out(2*NCALOFIFOS/2+5).eta,
                     merged_out_2_6_eta_V  => merged2_out(2*NCALOFIFOS/2+6).eta,
                     merged_out_2_7_eta_V  => merged2_out(2*NCALOFIFOS/2+7).eta,
                     merged_out_2_8_eta_V  => merged2_out(2*NCALOFIFOS/2+8).eta,
                     merged_out_2_9_eta_V  => merged2_out(2*NCALOFIFOS/2+9).eta,
                     merged_out_0_0_phi_V  => merged2_out(0*NCALOFIFOS/2+0).phi,
                     merged_out_0_1_phi_V  => merged2_out(0*NCALOFIFOS/2+1).phi,
                     merged_out_0_2_phi_V  => merged2_out(0*NCALOFIFOS/2+2).phi,
                     merged_out_0_3_phi_V  => merged2_out(0*NCALOFIFOS/2+3).phi,
                     merged_out_0_4_phi_V  => merged2_out(0*NCALOFIFOS/2+4).phi,
                     merged_out_0_5_phi_V  => merged2_out(0*NCALOFIFOS/2+5).phi,
                     merged_out_0_6_phi_V  => merged2_out(0*NCALOFIFOS/2+6).phi,
                     merged_out_0_7_phi_V  => merged2_out(0*NCALOFIFOS/2+7).phi,
                     merged_out_0_8_phi_V  => merged2_out(0*NCALOFIFOS/2+8).phi,
                     merged_out_0_9_phi_V  => merged2_out(0*NCALOFIFOS/2+9).phi,
                     merged_out_1_0_phi_V  => merged2_out(1*NCALOFIFOS/2+0).phi,
                     merged_out_1_1_phi_V  => merged2_out(1*NCALOFIFOS/2+1).phi,
                     merged_out_1_2_phi_V  => merged2_out(1*NCALOFIFOS/2+2).phi,
                     merged_out_1_3_phi_V  => merged2_out(1*NCALOFIFOS/2+3).phi,
                     merged_out_1_4_phi_V  => merged2_out(1*NCALOFIFOS/2+4).phi,
                     merged_out_1_5_phi_V  => merged2_out(1*NCALOFIFOS/2+5).phi,
                     merged_out_1_6_phi_V  => merged2_out(1*NCALOFIFOS/2+6).phi,
                     merged_out_1_7_phi_V  => merged2_out(1*NCALOFIFOS/2+7).phi,
                     merged_out_1_8_phi_V  => merged2_out(1*NCALOFIFOS/2+8).phi,
                     merged_out_1_9_phi_V  => merged2_out(1*NCALOFIFOS/2+9).phi,
                     merged_out_2_0_phi_V  => merged2_out(2*NCALOFIFOS/2+0).phi,
                     merged_out_2_1_phi_V  => merged2_out(2*NCALOFIFOS/2+1).phi,
                     merged_out_2_2_phi_V  => merged2_out(2*NCALOFIFOS/2+2).phi,
                     merged_out_2_3_phi_V  => merged2_out(2*NCALOFIFOS/2+3).phi,
                     merged_out_2_4_phi_V  => merged2_out(2*NCALOFIFOS/2+4).phi,
                     merged_out_2_5_phi_V  => merged2_out(2*NCALOFIFOS/2+5).phi,
                     merged_out_2_6_phi_V  => merged2_out(2*NCALOFIFOS/2+6).phi,
                     merged_out_2_7_phi_V  => merged2_out(2*NCALOFIFOS/2+7).phi,
                     merged_out_2_8_phi_V  => merged2_out(2*NCALOFIFOS/2+8).phi,
                     merged_out_2_9_phi_V  => merged2_out(2*NCALOFIFOS/2+9).phi,
                     merged_out_0_0_rest_V  => merged2_out(0*NCALOFIFOS/2+0).rest,
                     merged_out_0_1_rest_V  => merged2_out(0*NCALOFIFOS/2+1).rest,
                     merged_out_0_2_rest_V  => merged2_out(0*NCALOFIFOS/2+2).rest,
                     merged_out_0_3_rest_V  => merged2_out(0*NCALOFIFOS/2+3).rest,
                     merged_out_0_4_rest_V  => merged2_out(0*NCALOFIFOS/2+4).rest,
                     merged_out_0_5_rest_V  => merged2_out(0*NCALOFIFOS/2+5).rest,
                     merged_out_0_6_rest_V  => merged2_out(0*NCALOFIFOS/2+6).rest,
                     merged_out_0_7_rest_V  => merged2_out(0*NCALOFIFOS/2+7).rest,
                     merged_out_0_8_rest_V  => merged2_out(0*NCALOFIFOS/2+8).rest,
                     merged_out_0_9_rest_V  => merged2_out(0*NCALOFIFOS/2+9).rest,
                     merged_out_1_0_rest_V  => merged2_out(1*NCALOFIFOS/2+0).rest,
                     merged_out_1_1_rest_V  => merged2_out(1*NCALOFIFOS/2+1).rest,
                     merged_out_1_2_rest_V  => merged2_out(1*NCALOFIFOS/2+2).rest,
                     merged_out_1_3_rest_V  => merged2_out(1*NCALOFIFOS/2+3).rest,
                     merged_out_1_4_rest_V  => merged2_out(1*NCALOFIFOS/2+4).rest,
                     merged_out_1_5_rest_V  => merged2_out(1*NCALOFIFOS/2+5).rest,
                     merged_out_1_6_rest_V  => merged2_out(1*NCALOFIFOS/2+6).rest,
                     merged_out_1_7_rest_V  => merged2_out(1*NCALOFIFOS/2+7).rest,
                     merged_out_1_8_rest_V  => merged2_out(1*NCALOFIFOS/2+8).rest,
                     merged_out_1_9_rest_V  => merged2_out(1*NCALOFIFOS/2+9).rest,
                     merged_out_2_0_rest_V  => merged2_out(2*NCALOFIFOS/2+0).rest,
                     merged_out_2_1_rest_V  => merged2_out(2*NCALOFIFOS/2+1).rest,
                     merged_out_2_2_rest_V  => merged2_out(2*NCALOFIFOS/2+2).rest,
                     merged_out_2_3_rest_V  => merged2_out(2*NCALOFIFOS/2+3).rest,
                     merged_out_2_4_rest_V  => merged2_out(2*NCALOFIFOS/2+4).rest,
                     merged_out_2_5_rest_V  => merged2_out(2*NCALOFIFOS/2+5).rest,
                     merged_out_2_6_rest_V  => merged2_out(2*NCALOFIFOS/2+6).rest,
                     merged_out_2_7_rest_V  => merged2_out(2*NCALOFIFOS/2+7).rest,
                     merged_out_2_8_rest_V  => merged2_out(2*NCALOFIFOS/2+8).rest,
                     merged_out_2_9_rest_V  => merged2_out(2*NCALOFIFOS/2+9).rest,
                     merged_full_0_0  => merged2_full(0*NCALOFIFOS/2+0),
                     merged_full_0_1  => merged2_full(0*NCALOFIFOS/2+1),
                     merged_full_0_2  => merged2_full(0*NCALOFIFOS/2+2),
                     merged_full_0_3  => merged2_full(0*NCALOFIFOS/2+3),
                     merged_full_0_4  => merged2_full(0*NCALOFIFOS/2+4),
                     merged_full_0_5  => merged2_full(0*NCALOFIFOS/2+5),
                     merged_full_0_6  => merged2_full(0*NCALOFIFOS/2+6),
                     merged_full_0_7  => merged2_full(0*NCALOFIFOS/2+7),
                     merged_full_0_8  => merged2_full(0*NCALOFIFOS/2+8),
                     merged_full_0_9  => merged2_full(0*NCALOFIFOS/2+9),
                     merged_full_1_0  => merged2_full(1*NCALOFIFOS/2+0),
                     merged_full_1_1  => merged2_full(1*NCALOFIFOS/2+1),
                     merged_full_1_2  => merged2_full(1*NCALOFIFOS/2+2),
                     merged_full_1_3  => merged2_full(1*NCALOFIFOS/2+3),
                     merged_full_1_4  => merged2_full(1*NCALOFIFOS/2+4),
                     merged_full_1_5  => merged2_full(1*NCALOFIFOS/2+5),
                     merged_full_1_6  => merged2_full(1*NCALOFIFOS/2+6),
                     merged_full_1_7  => merged2_full(1*NCALOFIFOS/2+7),
                     merged_full_1_8  => merged2_full(1*NCALOFIFOS/2+8),
                     merged_full_1_9  => merged2_full(1*NCALOFIFOS/2+9),
                     merged_full_2_0  => merged2_full(2*NCALOFIFOS/2+0),
                     merged_full_2_1  => merged2_full(2*NCALOFIFOS/2+1),
                     merged_full_2_2  => merged2_full(2*NCALOFIFOS/2+2),
                     merged_full_2_3  => merged2_full(2*NCALOFIFOS/2+3),
                     merged_full_2_4  => merged2_full(2*NCALOFIFOS/2+4),
                     merged_full_2_5  => merged2_full(2*NCALOFIFOS/2+5),
                     merged_full_2_6  => merged2_full(2*NCALOFIFOS/2+6),
                     merged_full_2_7  => merged2_full(2*NCALOFIFOS/2+7),
                     merged_full_2_8  => merged2_full(2*NCALOFIFOS/2+8),
                     merged_full_2_9  => merged2_full(2*NCALOFIFOS/2+9),
                     merged_out_valid_0_0  => merged2_out_valid(0*NCALOFIFOS/2+0),
                     merged_out_valid_0_1  => merged2_out_valid(0*NCALOFIFOS/2+1),
                     merged_out_valid_0_2  => merged2_out_valid(0*NCALOFIFOS/2+2),
                     merged_out_valid_0_3  => merged2_out_valid(0*NCALOFIFOS/2+3),
                     merged_out_valid_0_4  => merged2_out_valid(0*NCALOFIFOS/2+4),
                     merged_out_valid_0_5  => merged2_out_valid(0*NCALOFIFOS/2+5),
                     merged_out_valid_0_6  => merged2_out_valid(0*NCALOFIFOS/2+6),
                     merged_out_valid_0_7  => merged2_out_valid(0*NCALOFIFOS/2+7),
                     merged_out_valid_0_8  => merged2_out_valid(0*NCALOFIFOS/2+8),
                     merged_out_valid_0_9  => merged2_out_valid(0*NCALOFIFOS/2+9),
                     merged_out_valid_1_0  => merged2_out_valid(1*NCALOFIFOS/2+0),
                     merged_out_valid_1_1  => merged2_out_valid(1*NCALOFIFOS/2+1),
                     merged_out_valid_1_2  => merged2_out_valid(1*NCALOFIFOS/2+2),
                     merged_out_valid_1_3  => merged2_out_valid(1*NCALOFIFOS/2+3),
                     merged_out_valid_1_4  => merged2_out_valid(1*NCALOFIFOS/2+4),
                     merged_out_valid_1_5  => merged2_out_valid(1*NCALOFIFOS/2+5),
                     merged_out_valid_1_6  => merged2_out_valid(1*NCALOFIFOS/2+6),
                     merged_out_valid_1_7  => merged2_out_valid(1*NCALOFIFOS/2+7),
                     merged_out_valid_1_8  => merged2_out_valid(1*NCALOFIFOS/2+8),
                     merged_out_valid_1_9  => merged2_out_valid(1*NCALOFIFOS/2+9),
                     merged_out_valid_2_0  => merged2_out_valid(2*NCALOFIFOS/2+0),
                     merged_out_valid_2_1  => merged2_out_valid(2*NCALOFIFOS/2+1),
                     merged_out_valid_2_2  => merged2_out_valid(2*NCALOFIFOS/2+2),
                     merged_out_valid_2_3  => merged2_out_valid(2*NCALOFIFOS/2+3),
                     merged_out_valid_2_4  => merged2_out_valid(2*NCALOFIFOS/2+4),
                     merged_out_valid_2_5  => merged2_out_valid(2*NCALOFIFOS/2+5),
                     merged_out_valid_2_6  => merged2_out_valid(2*NCALOFIFOS/2+6),
                     merged_out_valid_2_7  => merged2_out_valid(2*NCALOFIFOS/2+7),
                     merged_out_valid_2_8  => merged2_out_valid(2*NCALOFIFOS/2+8),
                     merged_out_valid_2_9  => merged2_out_valid(2*NCALOFIFOS/2+9),
                     merged_out_roll_0_0  => merged2_out_roll(0*NCALOFIFOS/2+0),
                     merged_out_roll_0_1  => merged2_out_roll(0*NCALOFIFOS/2+1),
                     merged_out_roll_0_2  => merged2_out_roll(0*NCALOFIFOS/2+2),
                     merged_out_roll_0_3  => merged2_out_roll(0*NCALOFIFOS/2+3),
                     merged_out_roll_0_4  => merged2_out_roll(0*NCALOFIFOS/2+4),
                     merged_out_roll_0_5  => merged2_out_roll(0*NCALOFIFOS/2+5),
                     merged_out_roll_0_6  => merged2_out_roll(0*NCALOFIFOS/2+6),
                     merged_out_roll_0_7  => merged2_out_roll(0*NCALOFIFOS/2+7),
                     merged_out_roll_0_8  => merged2_out_roll(0*NCALOFIFOS/2+8),
                     merged_out_roll_0_9  => merged2_out_roll(0*NCALOFIFOS/2+9),
                     merged_out_roll_1_0  => merged2_out_roll(1*NCALOFIFOS/2+0),
                     merged_out_roll_1_1  => merged2_out_roll(1*NCALOFIFOS/2+1),
                     merged_out_roll_1_2  => merged2_out_roll(1*NCALOFIFOS/2+2),
                     merged_out_roll_1_3  => merged2_out_roll(1*NCALOFIFOS/2+3),
                     merged_out_roll_1_4  => merged2_out_roll(1*NCALOFIFOS/2+4),
                     merged_out_roll_1_5  => merged2_out_roll(1*NCALOFIFOS/2+5),
                     merged_out_roll_1_6  => merged2_out_roll(1*NCALOFIFOS/2+6),
                     merged_out_roll_1_7  => merged2_out_roll(1*NCALOFIFOS/2+7),
                     merged_out_roll_1_8  => merged2_out_roll(1*NCALOFIFOS/2+8),
                     merged_out_roll_1_9  => merged2_out_roll(1*NCALOFIFOS/2+9),
                     merged_out_roll_2_0  => merged2_out_roll(2*NCALOFIFOS/2+0),
                     merged_out_roll_2_1  => merged2_out_roll(2*NCALOFIFOS/2+1),
                     merged_out_roll_2_2  => merged2_out_roll(2*NCALOFIFOS/2+2),
                     merged_out_roll_2_3  => merged2_out_roll(2*NCALOFIFOS/2+3),
                     merged_out_roll_2_4  => merged2_out_roll(2*NCALOFIFOS/2+4),
                     merged_out_roll_2_5  => merged2_out_roll(2*NCALOFIFOS/2+5),
                     merged_out_roll_2_6  => merged2_out_roll(2*NCALOFIFOS/2+6),
                     merged_out_roll_2_7  => merged2_out_roll(2*NCALOFIFOS/2+7),
                     merged_out_roll_2_8  => merged2_out_roll(2*NCALOFIFOS/2+8),
                     merged_out_roll_2_9  => merged2_out_roll(2*NCALOFIFOS/2+9)
                 );

  merge4_slice : entity work.calo_router_merge4_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     merged2_out_0_0_pt_V  => merged2_out(0*NCALOFIFOS/2+0).pt,
                     merged2_out_0_1_pt_V  => merged2_out(0*NCALOFIFOS/2+1).pt,
                     merged2_out_0_2_pt_V  => merged2_out(0*NCALOFIFOS/2+2).pt,
                     merged2_out_0_3_pt_V  => merged2_out(0*NCALOFIFOS/2+3).pt,
                     merged2_out_0_4_pt_V  => merged2_out(0*NCALOFIFOS/2+4).pt,
                     merged2_out_0_5_pt_V  => merged2_out(0*NCALOFIFOS/2+5).pt,
                     merged2_out_0_6_pt_V  => merged2_out(0*NCALOFIFOS/2+6).pt,
                     merged2_out_0_7_pt_V  => merged2_out(0*NCALOFIFOS/2+7).pt,
                     merged2_out_0_8_pt_V  => merged2_out(0*NCALOFIFOS/2+8).pt,
                     merged2_out_0_9_pt_V  => merged2_out(0*NCALOFIFOS/2+9).pt,
                     merged2_out_1_0_pt_V  => merged2_out(1*NCALOFIFOS/2+0).pt,
                     merged2_out_1_1_pt_V  => merged2_out(1*NCALOFIFOS/2+1).pt,
                     merged2_out_1_2_pt_V  => merged2_out(1*NCALOFIFOS/2+2).pt,
                     merged2_out_1_3_pt_V  => merged2_out(1*NCALOFIFOS/2+3).pt,
                     merged2_out_1_4_pt_V  => merged2_out(1*NCALOFIFOS/2+4).pt,
                     merged2_out_1_5_pt_V  => merged2_out(1*NCALOFIFOS/2+5).pt,
                     merged2_out_1_6_pt_V  => merged2_out(1*NCALOFIFOS/2+6).pt,
                     merged2_out_1_7_pt_V  => merged2_out(1*NCALOFIFOS/2+7).pt,
                     merged2_out_1_8_pt_V  => merged2_out(1*NCALOFIFOS/2+8).pt,
                     merged2_out_1_9_pt_V  => merged2_out(1*NCALOFIFOS/2+9).pt,
                     merged2_out_2_0_pt_V  => merged2_out(2*NCALOFIFOS/2+0).pt,
                     merged2_out_2_1_pt_V  => merged2_out(2*NCALOFIFOS/2+1).pt,
                     merged2_out_2_2_pt_V  => merged2_out(2*NCALOFIFOS/2+2).pt,
                     merged2_out_2_3_pt_V  => merged2_out(2*NCALOFIFOS/2+3).pt,
                     merged2_out_2_4_pt_V  => merged2_out(2*NCALOFIFOS/2+4).pt,
                     merged2_out_2_5_pt_V  => merged2_out(2*NCALOFIFOS/2+5).pt,
                     merged2_out_2_6_pt_V  => merged2_out(2*NCALOFIFOS/2+6).pt,
                     merged2_out_2_7_pt_V  => merged2_out(2*NCALOFIFOS/2+7).pt,
                     merged2_out_2_8_pt_V  => merged2_out(2*NCALOFIFOS/2+8).pt,
                     merged2_out_2_9_pt_V  => merged2_out(2*NCALOFIFOS/2+9).pt,
                     merged2_out_0_0_eta_V  => merged2_out(0*NCALOFIFOS/2+0).eta,
                     merged2_out_0_1_eta_V  => merged2_out(0*NCALOFIFOS/2+1).eta,
                     merged2_out_0_2_eta_V  => merged2_out(0*NCALOFIFOS/2+2).eta,
                     merged2_out_0_3_eta_V  => merged2_out(0*NCALOFIFOS/2+3).eta,
                     merged2_out_0_4_eta_V  => merged2_out(0*NCALOFIFOS/2+4).eta,
                     merged2_out_0_5_eta_V  => merged2_out(0*NCALOFIFOS/2+5).eta,
                     merged2_out_0_6_eta_V  => merged2_out(0*NCALOFIFOS/2+6).eta,
                     merged2_out_0_7_eta_V  => merged2_out(0*NCALOFIFOS/2+7).eta,
                     merged2_out_0_8_eta_V  => merged2_out(0*NCALOFIFOS/2+8).eta,
                     merged2_out_0_9_eta_V  => merged2_out(0*NCALOFIFOS/2+9).eta,
                     merged2_out_1_0_eta_V  => merged2_out(1*NCALOFIFOS/2+0).eta,
                     merged2_out_1_1_eta_V  => merged2_out(1*NCALOFIFOS/2+1).eta,
                     merged2_out_1_2_eta_V  => merged2_out(1*NCALOFIFOS/2+2).eta,
                     merged2_out_1_3_eta_V  => merged2_out(1*NCALOFIFOS/2+3).eta,
                     merged2_out_1_4_eta_V  => merged2_out(1*NCALOFIFOS/2+4).eta,
                     merged2_out_1_5_eta_V  => merged2_out(1*NCALOFIFOS/2+5).eta,
                     merged2_out_1_6_eta_V  => merged2_out(1*NCALOFIFOS/2+6).eta,
                     merged2_out_1_7_eta_V  => merged2_out(1*NCALOFIFOS/2+7).eta,
                     merged2_out_1_8_eta_V  => merged2_out(1*NCALOFIFOS/2+8).eta,
                     merged2_out_1_9_eta_V  => merged2_out(1*NCALOFIFOS/2+9).eta,
                     merged2_out_2_0_eta_V  => merged2_out(2*NCALOFIFOS/2+0).eta,
                     merged2_out_2_1_eta_V  => merged2_out(2*NCALOFIFOS/2+1).eta,
                     merged2_out_2_2_eta_V  => merged2_out(2*NCALOFIFOS/2+2).eta,
                     merged2_out_2_3_eta_V  => merged2_out(2*NCALOFIFOS/2+3).eta,
                     merged2_out_2_4_eta_V  => merged2_out(2*NCALOFIFOS/2+4).eta,
                     merged2_out_2_5_eta_V  => merged2_out(2*NCALOFIFOS/2+5).eta,
                     merged2_out_2_6_eta_V  => merged2_out(2*NCALOFIFOS/2+6).eta,
                     merged2_out_2_7_eta_V  => merged2_out(2*NCALOFIFOS/2+7).eta,
                     merged2_out_2_8_eta_V  => merged2_out(2*NCALOFIFOS/2+8).eta,
                     merged2_out_2_9_eta_V  => merged2_out(2*NCALOFIFOS/2+9).eta,
                     merged2_out_0_0_phi_V  => merged2_out(0*NCALOFIFOS/2+0).phi,
                     merged2_out_0_1_phi_V  => merged2_out(0*NCALOFIFOS/2+1).phi,
                     merged2_out_0_2_phi_V  => merged2_out(0*NCALOFIFOS/2+2).phi,
                     merged2_out_0_3_phi_V  => merged2_out(0*NCALOFIFOS/2+3).phi,
                     merged2_out_0_4_phi_V  => merged2_out(0*NCALOFIFOS/2+4).phi,
                     merged2_out_0_5_phi_V  => merged2_out(0*NCALOFIFOS/2+5).phi,
                     merged2_out_0_6_phi_V  => merged2_out(0*NCALOFIFOS/2+6).phi,
                     merged2_out_0_7_phi_V  => merged2_out(0*NCALOFIFOS/2+7).phi,
                     merged2_out_0_8_phi_V  => merged2_out(0*NCALOFIFOS/2+8).phi,
                     merged2_out_0_9_phi_V  => merged2_out(0*NCALOFIFOS/2+9).phi,
                     merged2_out_1_0_phi_V  => merged2_out(1*NCALOFIFOS/2+0).phi,
                     merged2_out_1_1_phi_V  => merged2_out(1*NCALOFIFOS/2+1).phi,
                     merged2_out_1_2_phi_V  => merged2_out(1*NCALOFIFOS/2+2).phi,
                     merged2_out_1_3_phi_V  => merged2_out(1*NCALOFIFOS/2+3).phi,
                     merged2_out_1_4_phi_V  => merged2_out(1*NCALOFIFOS/2+4).phi,
                     merged2_out_1_5_phi_V  => merged2_out(1*NCALOFIFOS/2+5).phi,
                     merged2_out_1_6_phi_V  => merged2_out(1*NCALOFIFOS/2+6).phi,
                     merged2_out_1_7_phi_V  => merged2_out(1*NCALOFIFOS/2+7).phi,
                     merged2_out_1_8_phi_V  => merged2_out(1*NCALOFIFOS/2+8).phi,
                     merged2_out_1_9_phi_V  => merged2_out(1*NCALOFIFOS/2+9).phi,
                     merged2_out_2_0_phi_V  => merged2_out(2*NCALOFIFOS/2+0).phi,
                     merged2_out_2_1_phi_V  => merged2_out(2*NCALOFIFOS/2+1).phi,
                     merged2_out_2_2_phi_V  => merged2_out(2*NCALOFIFOS/2+2).phi,
                     merged2_out_2_3_phi_V  => merged2_out(2*NCALOFIFOS/2+3).phi,
                     merged2_out_2_4_phi_V  => merged2_out(2*NCALOFIFOS/2+4).phi,
                     merged2_out_2_5_phi_V  => merged2_out(2*NCALOFIFOS/2+5).phi,
                     merged2_out_2_6_phi_V  => merged2_out(2*NCALOFIFOS/2+6).phi,
                     merged2_out_2_7_phi_V  => merged2_out(2*NCALOFIFOS/2+7).phi,
                     merged2_out_2_8_phi_V  => merged2_out(2*NCALOFIFOS/2+8).phi,
                     merged2_out_2_9_phi_V  => merged2_out(2*NCALOFIFOS/2+9).phi,
                     merged2_out_0_0_rest_V  => merged2_out(0*NCALOFIFOS/2+0).rest,
                     merged2_out_0_1_rest_V  => merged2_out(0*NCALOFIFOS/2+1).rest,
                     merged2_out_0_2_rest_V  => merged2_out(0*NCALOFIFOS/2+2).rest,
                     merged2_out_0_3_rest_V  => merged2_out(0*NCALOFIFOS/2+3).rest,
                     merged2_out_0_4_rest_V  => merged2_out(0*NCALOFIFOS/2+4).rest,
                     merged2_out_0_5_rest_V  => merged2_out(0*NCALOFIFOS/2+5).rest,
                     merged2_out_0_6_rest_V  => merged2_out(0*NCALOFIFOS/2+6).rest,
                     merged2_out_0_7_rest_V  => merged2_out(0*NCALOFIFOS/2+7).rest,
                     merged2_out_0_8_rest_V  => merged2_out(0*NCALOFIFOS/2+8).rest,
                     merged2_out_0_9_rest_V  => merged2_out(0*NCALOFIFOS/2+9).rest,
                     merged2_out_1_0_rest_V  => merged2_out(1*NCALOFIFOS/2+0).rest,
                     merged2_out_1_1_rest_V  => merged2_out(1*NCALOFIFOS/2+1).rest,
                     merged2_out_1_2_rest_V  => merged2_out(1*NCALOFIFOS/2+2).rest,
                     merged2_out_1_3_rest_V  => merged2_out(1*NCALOFIFOS/2+3).rest,
                     merged2_out_1_4_rest_V  => merged2_out(1*NCALOFIFOS/2+4).rest,
                     merged2_out_1_5_rest_V  => merged2_out(1*NCALOFIFOS/2+5).rest,
                     merged2_out_1_6_rest_V  => merged2_out(1*NCALOFIFOS/2+6).rest,
                     merged2_out_1_7_rest_V  => merged2_out(1*NCALOFIFOS/2+7).rest,
                     merged2_out_1_8_rest_V  => merged2_out(1*NCALOFIFOS/2+8).rest,
                     merged2_out_1_9_rest_V  => merged2_out(1*NCALOFIFOS/2+9).rest,
                     merged2_out_2_0_rest_V  => merged2_out(2*NCALOFIFOS/2+0).rest,
                     merged2_out_2_1_rest_V  => merged2_out(2*NCALOFIFOS/2+1).rest,
                     merged2_out_2_2_rest_V  => merged2_out(2*NCALOFIFOS/2+2).rest,
                     merged2_out_2_3_rest_V  => merged2_out(2*NCALOFIFOS/2+3).rest,
                     merged2_out_2_4_rest_V  => merged2_out(2*NCALOFIFOS/2+4).rest,
                     merged2_out_2_5_rest_V  => merged2_out(2*NCALOFIFOS/2+5).rest,
                     merged2_out_2_6_rest_V  => merged2_out(2*NCALOFIFOS/2+6).rest,
                     merged2_out_2_7_rest_V  => merged2_out(2*NCALOFIFOS/2+7).rest,
                     merged2_out_2_8_rest_V  => merged2_out(2*NCALOFIFOS/2+8).rest,
                     merged2_out_2_9_rest_V  => merged2_out(2*NCALOFIFOS/2+9).rest,
                     merged2_full_0_0  => merged2_full(0*NCALOFIFOS/2+0),
                     merged2_full_0_1  => merged2_full(0*NCALOFIFOS/2+1),
                     merged2_full_0_2  => merged2_full(0*NCALOFIFOS/2+2),
                     merged2_full_0_3  => merged2_full(0*NCALOFIFOS/2+3),
                     merged2_full_0_4  => merged2_full(0*NCALOFIFOS/2+4),
                     merged2_full_0_5  => merged2_full(0*NCALOFIFOS/2+5),
                     merged2_full_0_6  => merged2_full(0*NCALOFIFOS/2+6),
                     merged2_full_0_7  => merged2_full(0*NCALOFIFOS/2+7),
                     merged2_full_0_8  => merged2_full(0*NCALOFIFOS/2+8),
                     merged2_full_0_9  => merged2_full(0*NCALOFIFOS/2+9),
                     merged2_full_1_0  => merged2_full(1*NCALOFIFOS/2+0),
                     merged2_full_1_1  => merged2_full(1*NCALOFIFOS/2+1),
                     merged2_full_1_2  => merged2_full(1*NCALOFIFOS/2+2),
                     merged2_full_1_3  => merged2_full(1*NCALOFIFOS/2+3),
                     merged2_full_1_4  => merged2_full(1*NCALOFIFOS/2+4),
                     merged2_full_1_5  => merged2_full(1*NCALOFIFOS/2+5),
                     merged2_full_1_6  => merged2_full(1*NCALOFIFOS/2+6),
                     merged2_full_1_7  => merged2_full(1*NCALOFIFOS/2+7),
                     merged2_full_1_8  => merged2_full(1*NCALOFIFOS/2+8),
                     merged2_full_1_9  => merged2_full(1*NCALOFIFOS/2+9),
                     merged2_full_2_0  => merged2_full(2*NCALOFIFOS/2+0),
                     merged2_full_2_1  => merged2_full(2*NCALOFIFOS/2+1),
                     merged2_full_2_2  => merged2_full(2*NCALOFIFOS/2+2),
                     merged2_full_2_3  => merged2_full(2*NCALOFIFOS/2+3),
                     merged2_full_2_4  => merged2_full(2*NCALOFIFOS/2+4),
                     merged2_full_2_5  => merged2_full(2*NCALOFIFOS/2+5),
                     merged2_full_2_6  => merged2_full(2*NCALOFIFOS/2+6),
                     merged2_full_2_7  => merged2_full(2*NCALOFIFOS/2+7),
                     merged2_full_2_8  => merged2_full(2*NCALOFIFOS/2+8),
                     merged2_full_2_9  => merged2_full(2*NCALOFIFOS/2+9),
                     merged2_out_valid_0_0  => merged2_out_valid(0*NCALOFIFOS/2+0),
                     merged2_out_valid_0_1  => merged2_out_valid(0*NCALOFIFOS/2+1),
                     merged2_out_valid_0_2  => merged2_out_valid(0*NCALOFIFOS/2+2),
                     merged2_out_valid_0_3  => merged2_out_valid(0*NCALOFIFOS/2+3),
                     merged2_out_valid_0_4  => merged2_out_valid(0*NCALOFIFOS/2+4),
                     merged2_out_valid_0_5  => merged2_out_valid(0*NCALOFIFOS/2+5),
                     merged2_out_valid_0_6  => merged2_out_valid(0*NCALOFIFOS/2+6),
                     merged2_out_valid_0_7  => merged2_out_valid(0*NCALOFIFOS/2+7),
                     merged2_out_valid_0_8  => merged2_out_valid(0*NCALOFIFOS/2+8),
                     merged2_out_valid_0_9  => merged2_out_valid(0*NCALOFIFOS/2+9),
                     merged2_out_valid_1_0  => merged2_out_valid(1*NCALOFIFOS/2+0),
                     merged2_out_valid_1_1  => merged2_out_valid(1*NCALOFIFOS/2+1),
                     merged2_out_valid_1_2  => merged2_out_valid(1*NCALOFIFOS/2+2),
                     merged2_out_valid_1_3  => merged2_out_valid(1*NCALOFIFOS/2+3),
                     merged2_out_valid_1_4  => merged2_out_valid(1*NCALOFIFOS/2+4),
                     merged2_out_valid_1_5  => merged2_out_valid(1*NCALOFIFOS/2+5),
                     merged2_out_valid_1_6  => merged2_out_valid(1*NCALOFIFOS/2+6),
                     merged2_out_valid_1_7  => merged2_out_valid(1*NCALOFIFOS/2+7),
                     merged2_out_valid_1_8  => merged2_out_valid(1*NCALOFIFOS/2+8),
                     merged2_out_valid_1_9  => merged2_out_valid(1*NCALOFIFOS/2+9),
                     merged2_out_valid_2_0  => merged2_out_valid(2*NCALOFIFOS/2+0),
                     merged2_out_valid_2_1  => merged2_out_valid(2*NCALOFIFOS/2+1),
                     merged2_out_valid_2_2  => merged2_out_valid(2*NCALOFIFOS/2+2),
                     merged2_out_valid_2_3  => merged2_out_valid(2*NCALOFIFOS/2+3),
                     merged2_out_valid_2_4  => merged2_out_valid(2*NCALOFIFOS/2+4),
                     merged2_out_valid_2_5  => merged2_out_valid(2*NCALOFIFOS/2+5),
                     merged2_out_valid_2_6  => merged2_out_valid(2*NCALOFIFOS/2+6),
                     merged2_out_valid_2_7  => merged2_out_valid(2*NCALOFIFOS/2+7),
                     merged2_out_valid_2_8  => merged2_out_valid(2*NCALOFIFOS/2+8),
                     merged2_out_valid_2_9  => merged2_out_valid(2*NCALOFIFOS/2+9),
                     merged2_out_roll_0_0  => merged2_out_roll(0*NCALOFIFOS/2+0),
                     merged2_out_roll_0_1  => merged2_out_roll(0*NCALOFIFOS/2+1),
                     merged2_out_roll_0_2  => merged2_out_roll(0*NCALOFIFOS/2+2),
                     merged2_out_roll_0_3  => merged2_out_roll(0*NCALOFIFOS/2+3),
                     merged2_out_roll_0_4  => merged2_out_roll(0*NCALOFIFOS/2+4),
                     merged2_out_roll_0_5  => merged2_out_roll(0*NCALOFIFOS/2+5),
                     merged2_out_roll_0_6  => merged2_out_roll(0*NCALOFIFOS/2+6),
                     merged2_out_roll_0_7  => merged2_out_roll(0*NCALOFIFOS/2+7),
                     merged2_out_roll_0_8  => merged2_out_roll(0*NCALOFIFOS/2+8),
                     merged2_out_roll_0_9  => merged2_out_roll(0*NCALOFIFOS/2+9),
                     merged2_out_roll_1_0  => merged2_out_roll(1*NCALOFIFOS/2+0),
                     merged2_out_roll_1_1  => merged2_out_roll(1*NCALOFIFOS/2+1),
                     merged2_out_roll_1_2  => merged2_out_roll(1*NCALOFIFOS/2+2),
                     merged2_out_roll_1_3  => merged2_out_roll(1*NCALOFIFOS/2+3),
                     merged2_out_roll_1_4  => merged2_out_roll(1*NCALOFIFOS/2+4),
                     merged2_out_roll_1_5  => merged2_out_roll(1*NCALOFIFOS/2+5),
                     merged2_out_roll_1_6  => merged2_out_roll(1*NCALOFIFOS/2+6),
                     merged2_out_roll_1_7  => merged2_out_roll(1*NCALOFIFOS/2+7),
                     merged2_out_roll_1_8  => merged2_out_roll(1*NCALOFIFOS/2+8),
                     merged2_out_roll_1_9  => merged2_out_roll(1*NCALOFIFOS/2+9),
                     merged2_out_roll_2_0  => merged2_out_roll(2*NCALOFIFOS/2+0),
                     merged2_out_roll_2_1  => merged2_out_roll(2*NCALOFIFOS/2+1),
                     merged2_out_roll_2_2  => merged2_out_roll(2*NCALOFIFOS/2+2),
                     merged2_out_roll_2_3  => merged2_out_roll(2*NCALOFIFOS/2+3),
                     merged2_out_roll_2_4  => merged2_out_roll(2*NCALOFIFOS/2+4),
                     merged2_out_roll_2_5  => merged2_out_roll(2*NCALOFIFOS/2+5),
                     merged2_out_roll_2_6  => merged2_out_roll(2*NCALOFIFOS/2+6),
                     merged2_out_roll_2_7  => merged2_out_roll(2*NCALOFIFOS/2+7),
                     merged2_out_roll_2_8  => merged2_out_roll(2*NCALOFIFOS/2+8),
                     merged2_out_roll_2_9  => merged2_out_roll(2*NCALOFIFOS/2+9),
                     merged_out_0_0_pt_V  => merged4_out(0*NCALOFIFOS/4+0).pt,
                     merged_out_0_1_pt_V  => merged4_out(0*NCALOFIFOS/4+1).pt,
                     merged_out_0_2_pt_V  => merged4_out(0*NCALOFIFOS/4+2).pt,
                     merged_out_0_3_pt_V  => merged4_out(0*NCALOFIFOS/4+3).pt,
                     merged_out_0_4_pt_V  => merged4_out(0*NCALOFIFOS/4+4).pt,
                     merged_out_1_0_pt_V  => merged4_out(1*NCALOFIFOS/4+0).pt,
                     merged_out_1_1_pt_V  => merged4_out(1*NCALOFIFOS/4+1).pt,
                     merged_out_1_2_pt_V  => merged4_out(1*NCALOFIFOS/4+2).pt,
                     merged_out_1_3_pt_V  => merged4_out(1*NCALOFIFOS/4+3).pt,
                     merged_out_1_4_pt_V  => merged4_out(1*NCALOFIFOS/4+4).pt,
                     merged_out_2_0_pt_V  => merged4_out(2*NCALOFIFOS/4+0).pt,
                     merged_out_2_1_pt_V  => merged4_out(2*NCALOFIFOS/4+1).pt,
                     merged_out_2_2_pt_V  => merged4_out(2*NCALOFIFOS/4+2).pt,
                     merged_out_2_3_pt_V  => merged4_out(2*NCALOFIFOS/4+3).pt,
                     merged_out_2_4_pt_V  => merged4_out(2*NCALOFIFOS/4+4).pt,
                     merged_out_0_0_eta_V  => merged4_out(0*NCALOFIFOS/4+0).eta,
                     merged_out_0_1_eta_V  => merged4_out(0*NCALOFIFOS/4+1).eta,
                     merged_out_0_2_eta_V  => merged4_out(0*NCALOFIFOS/4+2).eta,
                     merged_out_0_3_eta_V  => merged4_out(0*NCALOFIFOS/4+3).eta,
                     merged_out_0_4_eta_V  => merged4_out(0*NCALOFIFOS/4+4).eta,
                     merged_out_1_0_eta_V  => merged4_out(1*NCALOFIFOS/4+0).eta,
                     merged_out_1_1_eta_V  => merged4_out(1*NCALOFIFOS/4+1).eta,
                     merged_out_1_2_eta_V  => merged4_out(1*NCALOFIFOS/4+2).eta,
                     merged_out_1_3_eta_V  => merged4_out(1*NCALOFIFOS/4+3).eta,
                     merged_out_1_4_eta_V  => merged4_out(1*NCALOFIFOS/4+4).eta,
                     merged_out_2_0_eta_V  => merged4_out(2*NCALOFIFOS/4+0).eta,
                     merged_out_2_1_eta_V  => merged4_out(2*NCALOFIFOS/4+1).eta,
                     merged_out_2_2_eta_V  => merged4_out(2*NCALOFIFOS/4+2).eta,
                     merged_out_2_3_eta_V  => merged4_out(2*NCALOFIFOS/4+3).eta,
                     merged_out_2_4_eta_V  => merged4_out(2*NCALOFIFOS/4+4).eta,
                     merged_out_0_0_phi_V  => merged4_out(0*NCALOFIFOS/4+0).phi,
                     merged_out_0_1_phi_V  => merged4_out(0*NCALOFIFOS/4+1).phi,
                     merged_out_0_2_phi_V  => merged4_out(0*NCALOFIFOS/4+2).phi,
                     merged_out_0_3_phi_V  => merged4_out(0*NCALOFIFOS/4+3).phi,
                     merged_out_0_4_phi_V  => merged4_out(0*NCALOFIFOS/4+4).phi,
                     merged_out_1_0_phi_V  => merged4_out(1*NCALOFIFOS/4+0).phi,
                     merged_out_1_1_phi_V  => merged4_out(1*NCALOFIFOS/4+1).phi,
                     merged_out_1_2_phi_V  => merged4_out(1*NCALOFIFOS/4+2).phi,
                     merged_out_1_3_phi_V  => merged4_out(1*NCALOFIFOS/4+3).phi,
                     merged_out_1_4_phi_V  => merged4_out(1*NCALOFIFOS/4+4).phi,
                     merged_out_2_0_phi_V  => merged4_out(2*NCALOFIFOS/4+0).phi,
                     merged_out_2_1_phi_V  => merged4_out(2*NCALOFIFOS/4+1).phi,
                     merged_out_2_2_phi_V  => merged4_out(2*NCALOFIFOS/4+2).phi,
                     merged_out_2_3_phi_V  => merged4_out(2*NCALOFIFOS/4+3).phi,
                     merged_out_2_4_phi_V  => merged4_out(2*NCALOFIFOS/4+4).phi,
                     merged_out_0_0_rest_V  => merged4_out(0*NCALOFIFOS/4+0).rest,
                     merged_out_0_1_rest_V  => merged4_out(0*NCALOFIFOS/4+1).rest,
                     merged_out_0_2_rest_V  => merged4_out(0*NCALOFIFOS/4+2).rest,
                     merged_out_0_3_rest_V  => merged4_out(0*NCALOFIFOS/4+3).rest,
                     merged_out_0_4_rest_V  => merged4_out(0*NCALOFIFOS/4+4).rest,
                     merged_out_1_0_rest_V  => merged4_out(1*NCALOFIFOS/4+0).rest,
                     merged_out_1_1_rest_V  => merged4_out(1*NCALOFIFOS/4+1).rest,
                     merged_out_1_2_rest_V  => merged4_out(1*NCALOFIFOS/4+2).rest,
                     merged_out_1_3_rest_V  => merged4_out(1*NCALOFIFOS/4+3).rest,
                     merged_out_1_4_rest_V  => merged4_out(1*NCALOFIFOS/4+4).rest,
                     merged_out_2_0_rest_V  => merged4_out(2*NCALOFIFOS/4+0).rest,
                     merged_out_2_1_rest_V  => merged4_out(2*NCALOFIFOS/4+1).rest,
                     merged_out_2_2_rest_V  => merged4_out(2*NCALOFIFOS/4+2).rest,
                     merged_out_2_3_rest_V  => merged4_out(2*NCALOFIFOS/4+3).rest,
                     merged_out_2_4_rest_V  => merged4_out(2*NCALOFIFOS/4+4).rest,
                     merged_full_0_0  => merged4_full(0*NCALOFIFOS/4+0),
                     merged_full_0_1  => merged4_full(0*NCALOFIFOS/4+1),
                     merged_full_0_2  => merged4_full(0*NCALOFIFOS/4+2),
                     merged_full_0_3  => merged4_full(0*NCALOFIFOS/4+3),
                     merged_full_0_4  => merged4_full(0*NCALOFIFOS/4+4),
                     merged_full_1_0  => merged4_full(1*NCALOFIFOS/4+0),
                     merged_full_1_1  => merged4_full(1*NCALOFIFOS/4+1),
                     merged_full_1_2  => merged4_full(1*NCALOFIFOS/4+2),
                     merged_full_1_3  => merged4_full(1*NCALOFIFOS/4+3),
                     merged_full_1_4  => merged4_full(1*NCALOFIFOS/4+4),
                     merged_full_2_0  => merged4_full(2*NCALOFIFOS/4+0),
                     merged_full_2_1  => merged4_full(2*NCALOFIFOS/4+1),
                     merged_full_2_2  => merged4_full(2*NCALOFIFOS/4+2),
                     merged_full_2_3  => merged4_full(2*NCALOFIFOS/4+3),
                     merged_full_2_4  => merged4_full(2*NCALOFIFOS/4+4),
                     merged_out_valid_0_0  => merged4_out_valid(0*NCALOFIFOS/4+0),
                     merged_out_valid_0_1  => merged4_out_valid(0*NCALOFIFOS/4+1),
                     merged_out_valid_0_2  => merged4_out_valid(0*NCALOFIFOS/4+2),
                     merged_out_valid_0_3  => merged4_out_valid(0*NCALOFIFOS/4+3),
                     merged_out_valid_0_4  => merged4_out_valid(0*NCALOFIFOS/4+4),
                     merged_out_valid_1_0  => merged4_out_valid(1*NCALOFIFOS/4+0),
                     merged_out_valid_1_1  => merged4_out_valid(1*NCALOFIFOS/4+1),
                     merged_out_valid_1_2  => merged4_out_valid(1*NCALOFIFOS/4+2),
                     merged_out_valid_1_3  => merged4_out_valid(1*NCALOFIFOS/4+3),
                     merged_out_valid_1_4  => merged4_out_valid(1*NCALOFIFOS/4+4),
                     merged_out_valid_2_0  => merged4_out_valid(2*NCALOFIFOS/4+0),
                     merged_out_valid_2_1  => merged4_out_valid(2*NCALOFIFOS/4+1),
                     merged_out_valid_2_2  => merged4_out_valid(2*NCALOFIFOS/4+2),
                     merged_out_valid_2_3  => merged4_out_valid(2*NCALOFIFOS/4+3),
                     merged_out_valid_2_4  => merged4_out_valid(2*NCALOFIFOS/4+4),
                     merged_out_roll_0_0  => merged4_out_roll(0*NCALOFIFOS/4+0),
                     merged_out_roll_0_1  => merged4_out_roll(0*NCALOFIFOS/4+1),
                     merged_out_roll_0_2  => merged4_out_roll(0*NCALOFIFOS/4+2),
                     merged_out_roll_0_3  => merged4_out_roll(0*NCALOFIFOS/4+3),
                     merged_out_roll_0_4  => merged4_out_roll(0*NCALOFIFOS/4+4),
                     merged_out_roll_1_0  => merged4_out_roll(1*NCALOFIFOS/4+0),
                     merged_out_roll_1_1  => merged4_out_roll(1*NCALOFIFOS/4+1),
                     merged_out_roll_1_2  => merged4_out_roll(1*NCALOFIFOS/4+2),
                     merged_out_roll_1_3  => merged4_out_roll(1*NCALOFIFOS/4+3),
                     merged_out_roll_1_4  => merged4_out_roll(1*NCALOFIFOS/4+4),
                     merged_out_roll_2_0  => merged4_out_roll(2*NCALOFIFOS/4+0),
                     merged_out_roll_2_1  => merged4_out_roll(2*NCALOFIFOS/4+1),
                     merged_out_roll_2_2  => merged4_out_roll(2*NCALOFIFOS/4+2),
                     merged_out_roll_2_3  => merged4_out_roll(2*NCALOFIFOS/4+3),
                     merged_out_roll_2_4  => merged4_out_roll(2*NCALOFIFOS/4+4)
             );

            
            
  merge_slice : entity work.calo_router_merge_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     merged4_out_0_0_pt_V  => merged4_out(0*NCALOFIFOS/4+0).pt,
                     merged4_out_0_1_pt_V  => merged4_out(0*NCALOFIFOS/4+1).pt,
                     merged4_out_0_2_pt_V  => merged4_out(0*NCALOFIFOS/4+2).pt,
                     merged4_out_0_3_pt_V  => merged4_out(0*NCALOFIFOS/4+3).pt,
                     merged4_out_0_4_pt_V  => merged4_out(0*NCALOFIFOS/4+4).pt,
                     merged4_out_1_0_pt_V  => merged4_out(1*NCALOFIFOS/4+0).pt,
                     merged4_out_1_1_pt_V  => merged4_out(1*NCALOFIFOS/4+1).pt,
                     merged4_out_1_2_pt_V  => merged4_out(1*NCALOFIFOS/4+2).pt,
                     merged4_out_1_3_pt_V  => merged4_out(1*NCALOFIFOS/4+3).pt,
                     merged4_out_1_4_pt_V  => merged4_out(1*NCALOFIFOS/4+4).pt,
                     merged4_out_2_0_pt_V  => merged4_out(2*NCALOFIFOS/4+0).pt,
                     merged4_out_2_1_pt_V  => merged4_out(2*NCALOFIFOS/4+1).pt,
                     merged4_out_2_2_pt_V  => merged4_out(2*NCALOFIFOS/4+2).pt,
                     merged4_out_2_3_pt_V  => merged4_out(2*NCALOFIFOS/4+3).pt,
                     merged4_out_2_4_pt_V  => merged4_out(2*NCALOFIFOS/4+4).pt,
                     merged4_out_0_0_eta_V  => merged4_out(0*NCALOFIFOS/4+0).eta,
                     merged4_out_0_1_eta_V  => merged4_out(0*NCALOFIFOS/4+1).eta,
                     merged4_out_0_2_eta_V  => merged4_out(0*NCALOFIFOS/4+2).eta,
                     merged4_out_0_3_eta_V  => merged4_out(0*NCALOFIFOS/4+3).eta,
                     merged4_out_0_4_eta_V  => merged4_out(0*NCALOFIFOS/4+4).eta,
                     merged4_out_1_0_eta_V  => merged4_out(1*NCALOFIFOS/4+0).eta,
                     merged4_out_1_1_eta_V  => merged4_out(1*NCALOFIFOS/4+1).eta,
                     merged4_out_1_2_eta_V  => merged4_out(1*NCALOFIFOS/4+2).eta,
                     merged4_out_1_3_eta_V  => merged4_out(1*NCALOFIFOS/4+3).eta,
                     merged4_out_1_4_eta_V  => merged4_out(1*NCALOFIFOS/4+4).eta,
                     merged4_out_2_0_eta_V  => merged4_out(2*NCALOFIFOS/4+0).eta,
                     merged4_out_2_1_eta_V  => merged4_out(2*NCALOFIFOS/4+1).eta,
                     merged4_out_2_2_eta_V  => merged4_out(2*NCALOFIFOS/4+2).eta,
                     merged4_out_2_3_eta_V  => merged4_out(2*NCALOFIFOS/4+3).eta,
                     merged4_out_2_4_eta_V  => merged4_out(2*NCALOFIFOS/4+4).eta,
                     merged4_out_0_0_phi_V  => merged4_out(0*NCALOFIFOS/4+0).phi,
                     merged4_out_0_1_phi_V  => merged4_out(0*NCALOFIFOS/4+1).phi,
                     merged4_out_0_2_phi_V  => merged4_out(0*NCALOFIFOS/4+2).phi,
                     merged4_out_0_3_phi_V  => merged4_out(0*NCALOFIFOS/4+3).phi,
                     merged4_out_0_4_phi_V  => merged4_out(0*NCALOFIFOS/4+4).phi,
                     merged4_out_1_0_phi_V  => merged4_out(1*NCALOFIFOS/4+0).phi,
                     merged4_out_1_1_phi_V  => merged4_out(1*NCALOFIFOS/4+1).phi,
                     merged4_out_1_2_phi_V  => merged4_out(1*NCALOFIFOS/4+2).phi,
                     merged4_out_1_3_phi_V  => merged4_out(1*NCALOFIFOS/4+3).phi,
                     merged4_out_1_4_phi_V  => merged4_out(1*NCALOFIFOS/4+4).phi,
                     merged4_out_2_0_phi_V  => merged4_out(2*NCALOFIFOS/4+0).phi,
                     merged4_out_2_1_phi_V  => merged4_out(2*NCALOFIFOS/4+1).phi,
                     merged4_out_2_2_phi_V  => merged4_out(2*NCALOFIFOS/4+2).phi,
                     merged4_out_2_3_phi_V  => merged4_out(2*NCALOFIFOS/4+3).phi,
                     merged4_out_2_4_phi_V  => merged4_out(2*NCALOFIFOS/4+4).phi,
                     merged4_out_0_0_rest_V  => merged4_out(0*NCALOFIFOS/4+0).rest,
                     merged4_out_0_1_rest_V  => merged4_out(0*NCALOFIFOS/4+1).rest,
                     merged4_out_0_2_rest_V  => merged4_out(0*NCALOFIFOS/4+2).rest,
                     merged4_out_0_3_rest_V  => merged4_out(0*NCALOFIFOS/4+3).rest,
                     merged4_out_0_4_rest_V  => merged4_out(0*NCALOFIFOS/4+4).rest,
                     merged4_out_1_0_rest_V  => merged4_out(1*NCALOFIFOS/4+0).rest,
                     merged4_out_1_1_rest_V  => merged4_out(1*NCALOFIFOS/4+1).rest,
                     merged4_out_1_2_rest_V  => merged4_out(1*NCALOFIFOS/4+2).rest,
                     merged4_out_1_3_rest_V  => merged4_out(1*NCALOFIFOS/4+3).rest,
                     merged4_out_1_4_rest_V  => merged4_out(1*NCALOFIFOS/4+4).rest,
                     merged4_out_2_0_rest_V  => merged4_out(2*NCALOFIFOS/4+0).rest,
                     merged4_out_2_1_rest_V  => merged4_out(2*NCALOFIFOS/4+1).rest,
                     merged4_out_2_2_rest_V  => merged4_out(2*NCALOFIFOS/4+2).rest,
                     merged4_out_2_3_rest_V  => merged4_out(2*NCALOFIFOS/4+3).rest,
                     merged4_out_2_4_rest_V  => merged4_out(2*NCALOFIFOS/4+4).rest,
                     merged4_full_0_0  => merged4_full(0*NCALOFIFOS/4+0),
                     merged4_full_0_1  => merged4_full(0*NCALOFIFOS/4+1),
                     merged4_full_0_2  => merged4_full(0*NCALOFIFOS/4+2),
                     merged4_full_0_3  => merged4_full(0*NCALOFIFOS/4+3),
                     merged4_full_0_4  => merged4_full(0*NCALOFIFOS/4+4),
                     merged4_full_1_0  => merged4_full(1*NCALOFIFOS/4+0),
                     merged4_full_1_1  => merged4_full(1*NCALOFIFOS/4+1),
                     merged4_full_1_2  => merged4_full(1*NCALOFIFOS/4+2),
                     merged4_full_1_3  => merged4_full(1*NCALOFIFOS/4+3),
                     merged4_full_1_4  => merged4_full(1*NCALOFIFOS/4+4),
                     merged4_full_2_0  => merged4_full(2*NCALOFIFOS/4+0),
                     merged4_full_2_1  => merged4_full(2*NCALOFIFOS/4+1),
                     merged4_full_2_2  => merged4_full(2*NCALOFIFOS/4+2),
                     merged4_full_2_3  => merged4_full(2*NCALOFIFOS/4+3),
                     merged4_full_2_4  => merged4_full(2*NCALOFIFOS/4+4),
                     merged4_out_valid_0_0  => merged4_out_valid(0*NCALOFIFOS/4+0),
                     merged4_out_valid_0_1  => merged4_out_valid(0*NCALOFIFOS/4+1),
                     merged4_out_valid_0_2  => merged4_out_valid(0*NCALOFIFOS/4+2),
                     merged4_out_valid_0_3  => merged4_out_valid(0*NCALOFIFOS/4+3),
                     merged4_out_valid_0_4  => merged4_out_valid(0*NCALOFIFOS/4+4),
                     merged4_out_valid_1_0  => merged4_out_valid(1*NCALOFIFOS/4+0),
                     merged4_out_valid_1_1  => merged4_out_valid(1*NCALOFIFOS/4+1),
                     merged4_out_valid_1_2  => merged4_out_valid(1*NCALOFIFOS/4+2),
                     merged4_out_valid_1_3  => merged4_out_valid(1*NCALOFIFOS/4+3),
                     merged4_out_valid_1_4  => merged4_out_valid(1*NCALOFIFOS/4+4),
                     merged4_out_valid_2_0  => merged4_out_valid(2*NCALOFIFOS/4+0),
                     merged4_out_valid_2_1  => merged4_out_valid(2*NCALOFIFOS/4+1),
                     merged4_out_valid_2_2  => merged4_out_valid(2*NCALOFIFOS/4+2),
                     merged4_out_valid_2_3  => merged4_out_valid(2*NCALOFIFOS/4+3),
                     merged4_out_valid_2_4  => merged4_out_valid(2*NCALOFIFOS/4+4),
                     merged4_out_roll_0_0  => merged4_out_roll(0*NCALOFIFOS/4+0),
                     merged4_out_roll_0_1  => merged4_out_roll(0*NCALOFIFOS/4+1),
                     merged4_out_roll_0_2  => merged4_out_roll(0*NCALOFIFOS/4+2),
                     merged4_out_roll_0_3  => merged4_out_roll(0*NCALOFIFOS/4+3),
                     merged4_out_roll_0_4  => merged4_out_roll(0*NCALOFIFOS/4+4),
                     merged4_out_roll_1_0  => merged4_out_roll(1*NCALOFIFOS/4+0),
                     merged4_out_roll_1_1  => merged4_out_roll(1*NCALOFIFOS/4+1),
                     merged4_out_roll_1_2  => merged4_out_roll(1*NCALOFIFOS/4+2),
                     merged4_out_roll_1_3  => merged4_out_roll(1*NCALOFIFOS/4+3),
                     merged4_out_roll_1_4  => merged4_out_roll(1*NCALOFIFOS/4+4),
                     merged4_out_roll_2_0  => merged4_out_roll(2*NCALOFIFOS/4+0),
                     merged4_out_roll_2_1  => merged4_out_roll(2*NCALOFIFOS/4+1),
                     merged4_out_roll_2_2  => merged4_out_roll(2*NCALOFIFOS/4+2),
                     merged4_out_roll_2_3  => merged4_out_roll(2*NCALOFIFOS/4+3),
                     merged4_out_roll_2_4  => merged4_out_roll(2*NCALOFIFOS/4+4),
                     merged_out_0_pt_V  => merged_out(0).pt,
                     merged_out_1_pt_V  => merged_out(1).pt,
                     merged_out_2_pt_V  => merged_out(2).pt,
                     merged_out_3_pt_V  => merged_out(3).pt,
                     merged_out_4_pt_V  => merged_out(4).pt,
                     merged_out_5_pt_V  => merged_out(5).pt,
                     merged_out_6_pt_V  => merged_out(6).pt,
                     merged_out_7_pt_V  => merged_out(7).pt,
                     merged_out_8_pt_V  => merged_out(8).pt,
                     merged_out_0_eta_V  => merged_out(0).eta,
                     merged_out_1_eta_V  => merged_out(1).eta,
                     merged_out_2_eta_V  => merged_out(2).eta,
                     merged_out_3_eta_V  => merged_out(3).eta,
                     merged_out_4_eta_V  => merged_out(4).eta,
                     merged_out_5_eta_V  => merged_out(5).eta,
                     merged_out_6_eta_V  => merged_out(6).eta,
                     merged_out_7_eta_V  => merged_out(7).eta,
                     merged_out_8_eta_V  => merged_out(8).eta,
                     merged_out_0_phi_V  => merged_out(0).phi,
                     merged_out_1_phi_V  => merged_out(1).phi,
                     merged_out_2_phi_V  => merged_out(2).phi,
                     merged_out_3_phi_V  => merged_out(3).phi,
                     merged_out_4_phi_V  => merged_out(4).phi,
                     merged_out_5_phi_V  => merged_out(5).phi,
                     merged_out_6_phi_V  => merged_out(6).phi,
                     merged_out_7_phi_V  => merged_out(7).phi,
                     merged_out_8_phi_V  => merged_out(8).phi,
                     merged_out_0_rest_V  => merged_out(0).rest,
                     merged_out_1_rest_V  => merged_out(1).rest,
                     merged_out_2_rest_V  => merged_out(2).rest,
                     merged_out_3_rest_V  => merged_out(3).rest,
                     merged_out_4_rest_V  => merged_out(4).rest,
                     merged_out_5_rest_V  => merged_out(5).rest,
                     merged_out_6_rest_V  => merged_out(6).rest,
                     merged_out_7_rest_V  => merged_out(7).rest,
                     merged_out_8_rest_V  => merged_out(8).rest,
                     merged_out_valid_0  => merged_out_valid(0),
                     merged_out_valid_1  => merged_out_valid(1),
                     merged_out_valid_2  => merged_out_valid(2),
                     merged_out_valid_3  => merged_out_valid(3),
                     merged_out_valid_4  => merged_out_valid(4),
                     merged_out_valid_5  => merged_out_valid(5),
                     merged_out_valid_6  => merged_out_valid(6),
                     merged_out_valid_7  => merged_out_valid(7),
                     merged_out_valid_8  => merged_out_valid(8),
                     merged_out_roll_0  => merged_out_roll(0),
                     merged_out_roll_1  => merged_out_roll(1),
                     merged_out_roll_2  => merged_out_roll(2),
                     merged_out_roll_3  => merged_out_roll(3),
                     merged_out_roll_4  => merged_out_roll(4),
                     merged_out_roll_5  => merged_out_roll(5),
                     merged_out_roll_6  => merged_out_roll(6),
                     merged_out_roll_7  => merged_out_roll(7),
                     merged_out_roll_8  => merged_out_roll(8)
                );

  output_slice : entity work.calo_router_full_output_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     merged_out_0_pt_V  => merged_out(0).pt,
                     merged_out_1_pt_V  => merged_out(1).pt,
                     merged_out_2_pt_V  => merged_out(2).pt,
                     merged_out_3_pt_V  => merged_out(3).pt,
                     merged_out_4_pt_V  => merged_out(4).pt,
                     merged_out_5_pt_V  => merged_out(5).pt,
                     merged_out_6_pt_V  => merged_out(6).pt,
                     merged_out_7_pt_V  => merged_out(7).pt,
                     merged_out_8_pt_V  => merged_out(8).pt,
                     merged_out_0_eta_V  => merged_out(0).eta,
                     merged_out_1_eta_V  => merged_out(1).eta,
                     merged_out_2_eta_V  => merged_out(2).eta,
                     merged_out_3_eta_V  => merged_out(3).eta,
                     merged_out_4_eta_V  => merged_out(4).eta,
                     merged_out_5_eta_V  => merged_out(5).eta,
                     merged_out_6_eta_V  => merged_out(6).eta,
                     merged_out_7_eta_V  => merged_out(7).eta,
                     merged_out_8_eta_V  => merged_out(8).eta,
                     merged_out_0_phi_V  => merged_out(0).phi,
                     merged_out_1_phi_V  => merged_out(1).phi,
                     merged_out_2_phi_V  => merged_out(2).phi,
                     merged_out_3_phi_V  => merged_out(3).phi,
                     merged_out_4_phi_V  => merged_out(4).phi,
                     merged_out_5_phi_V  => merged_out(5).phi,
                     merged_out_6_phi_V  => merged_out(6).phi,
                     merged_out_7_phi_V  => merged_out(7).phi,
                     merged_out_8_phi_V  => merged_out(8).phi,
                     merged_out_0_rest_V  => merged_out(0).rest,
                     merged_out_1_rest_V  => merged_out(1).rest,
                     merged_out_2_rest_V  => merged_out(2).rest,
                     merged_out_3_rest_V  => merged_out(3).rest,
                     merged_out_4_rest_V  => merged_out(4).rest,
                     merged_out_5_rest_V  => merged_out(5).rest,
                     merged_out_6_rest_V  => merged_out(6).rest,
                     merged_out_7_rest_V  => merged_out(7).rest,
                     merged_out_8_rest_V  => merged_out(8).rest,
                     merged_out_valid_0  => merged_out_valid(0),
                     merged_out_valid_1  => merged_out_valid(1),
                     merged_out_valid_2  => merged_out_valid(2),
                     merged_out_valid_3  => merged_out_valid(3),
                     merged_out_valid_4  => merged_out_valid(4),
                     merged_out_valid_5  => merged_out_valid(5),
                     merged_out_valid_6  => merged_out_valid(6),
                     merged_out_valid_7  => merged_out_valid(7),
                     merged_out_valid_8  => merged_out_valid(8),
                     merged_out_roll_0  => merged_out_roll(0),
                     merged_out_roll_1  => merged_out_roll(1),
                     merged_out_roll_2  => merged_out_roll(2),
                     merged_out_roll_3  => merged_out_roll(3),
                     merged_out_roll_4  => merged_out_roll(4),
                     merged_out_roll_5  => merged_out_roll(5),
                     merged_out_roll_6  => merged_out_roll(6),
                     merged_out_roll_7  => merged_out_roll(7),
                     merged_out_roll_8  => merged_out_roll(8),
                     tracks_out_0_pt_V => tracks_out_0_pt_V,
                     tracks_out_1_pt_V => tracks_out_1_pt_V,
                     tracks_out_2_pt_V => tracks_out_2_pt_V,
                     tracks_out_3_pt_V => tracks_out_3_pt_V,
                     tracks_out_4_pt_V => tracks_out_4_pt_V,
                     tracks_out_5_pt_V => tracks_out_5_pt_V,
                     tracks_out_6_pt_V => tracks_out_6_pt_V,
                     tracks_out_7_pt_V => tracks_out_7_pt_V,
                     tracks_out_8_pt_V => tracks_out_8_pt_V,
                     tracks_out_0_eta_V => tracks_out_0_eta_V,
                     tracks_out_1_eta_V => tracks_out_1_eta_V,
                     tracks_out_2_eta_V => tracks_out_2_eta_V,
                     tracks_out_3_eta_V => tracks_out_3_eta_V,
                     tracks_out_4_eta_V => tracks_out_4_eta_V,
                     tracks_out_5_eta_V => tracks_out_5_eta_V,
                     tracks_out_6_eta_V => tracks_out_6_eta_V,
                     tracks_out_7_eta_V => tracks_out_7_eta_V,
                     tracks_out_8_eta_V => tracks_out_8_eta_V,
                     tracks_out_0_phi_V => tracks_out_0_phi_V,
                     tracks_out_1_phi_V => tracks_out_1_phi_V,
                     tracks_out_2_phi_V => tracks_out_2_phi_V,
                     tracks_out_3_phi_V => tracks_out_3_phi_V,
                     tracks_out_4_phi_V => tracks_out_4_phi_V,
                     tracks_out_5_phi_V => tracks_out_5_phi_V,
                     tracks_out_6_phi_V => tracks_out_6_phi_V,
                     tracks_out_7_phi_V => tracks_out_7_phi_V,
                     tracks_out_8_phi_V => tracks_out_8_phi_V,
                     tracks_out_0_rest_V => tracks_out_0_rest_V,
                     tracks_out_1_rest_V => tracks_out_1_rest_V,
                     tracks_out_2_rest_V => tracks_out_2_rest_V,
                     tracks_out_3_rest_V => tracks_out_3_rest_V,
                     tracks_out_4_rest_V => tracks_out_4_rest_V,
                     tracks_out_5_rest_V => tracks_out_5_rest_V,
                     tracks_out_6_rest_V => tracks_out_6_rest_V,
                     tracks_out_7_rest_V => tracks_out_7_rest_V,
                     tracks_out_8_rest_V => tracks_out_8_rest_V,
                     newevent_out => newevent_out
                );
end Behavioral;
