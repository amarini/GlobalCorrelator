library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.regionizer_data.all;

entity regionizer is
    port(
            ap_clk : IN STD_LOGIC;
            ap_rst : IN STD_LOGIC;
            ap_start : IN STD_LOGIC;
            ap_done : OUT STD_LOGIC;
            ap_idle : OUT STD_LOGIC;
            ap_ready : OUT STD_LOGIC;
            newevent : IN STD_LOGIC;
            tracks_in_0_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_1_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_2_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_0_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_1_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_2_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_0_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_0_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_1_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_2_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_3_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_3_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_4_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_4_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_5_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_5_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_3_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_4_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_5_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_3_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_3_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_4_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_4_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_5_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_5_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_6_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_6_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_7_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_7_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_8_0_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_8_1_pt_V : IN STD_LOGIC_VECTOR (13 downto 0);
            tracks_in_6_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_0_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_1_eta_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_7_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_0_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_8_1_phi_V : IN STD_LOGIC_VECTOR (11 downto 0);
            tracks_in_6_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_6_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_7_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_7_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_8_0_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_in_8_1_rest_V : IN STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_0_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_0_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_0_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_1_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_1_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_1_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_2_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_2_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_2_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_3_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_3_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_3_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_4_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_4_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_4_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_5_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_5_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_5_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_6_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_6_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_6_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_7_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_7_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_7_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            tracks_out_8_eta_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_phi_V : OUT STD_LOGIC_VECTOR (11 downto 0);
            tracks_out_8_pt_V : OUT STD_LOGIC_VECTOR (13 downto 0);
            tracks_out_8_rest_V : OUT STD_LOGIC_VECTOR (25 downto 0);
            newevent_out : OUT STD_LOGIC

    );
end regionizer;

architecture Behavioral of regionizer is
    constant NMERGED2  : natural := NSECTORS*(NFIFOS/2);
    constant NALLFIFOS : natural := NSECTORS*NFIFOS;
    constant NREGIONS  : natural := NSECTORS;

    signal links_in :       particles(NSECTORS*NFIBERS-1 downto 0);
    signal fifo_in :        particles(NALLFIFOS-1 downto 0);
    signal fifo_in_write :  std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');
    signal fifo_in_roll  :  std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');

    signal fifo_out :         particles(NALLFIFOS-1 downto 0);
    signal fifo_out_valid :   std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');
    signal fifo_out_full:     std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');
    signal fifo_out_roll:     std_logic_vector(NALLFIFOS-1 downto 0) := (others => '0');

    signal merged2_out :        particles(NMERGED2-1 downto 0);
    signal merged2_out_valid :  std_logic_vector(NMERGED2-1 downto 0) := (others => '0');
    signal merged2_out_roll:    std_logic_vector(NMERGED2-1 downto 0) := (others => '0');
    signal merged2_full:        std_logic_vector(NMERGED2-1 downto 0) := (others => '0');

    signal merged_out :        particles(NREGIONS-1 downto 0);
    signal merged_out_valid :  std_logic_vector(NREGIONS-1 downto 0) := (others => '0');
    signal merged_out_roll:    std_logic_vector(NREGIONS-1 downto 0) := (others => '0');

    signal newevent_del : std_logic;
begin

    delay : process (ap_clk)
    begin
        if rising_edge(ap_clk) then
            newevent_del <= newevent;
        end if;
    end process delay;

    input_slice : entity work.router_input_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     tracks_in_0_0_pt_V => tracks_in_0_0_pt_V,
                     tracks_in_0_1_pt_V => tracks_in_0_1_pt_V,
                     tracks_in_1_0_pt_V => tracks_in_1_0_pt_V,
                     tracks_in_1_1_pt_V => tracks_in_1_1_pt_V,
                     tracks_in_2_0_pt_V => tracks_in_2_0_pt_V,
                     tracks_in_2_1_pt_V => tracks_in_2_1_pt_V,
                     tracks_in_3_0_pt_V => tracks_in_3_0_pt_V,
                     tracks_in_3_1_pt_V => tracks_in_3_1_pt_V,
                     tracks_in_4_0_pt_V => tracks_in_4_0_pt_V,
                     tracks_in_4_1_pt_V => tracks_in_4_1_pt_V,
                     tracks_in_5_0_pt_V => tracks_in_5_0_pt_V,
                     tracks_in_5_1_pt_V => tracks_in_5_1_pt_V,
                     tracks_in_6_0_pt_V => tracks_in_6_0_pt_V,
                     tracks_in_6_1_pt_V => tracks_in_6_1_pt_V,
                     tracks_in_7_0_pt_V => tracks_in_7_0_pt_V,
                     tracks_in_7_1_pt_V => tracks_in_7_1_pt_V,
                     tracks_in_8_0_pt_V => tracks_in_8_0_pt_V,
                     tracks_in_8_1_pt_V => tracks_in_8_1_pt_V,
                     tracks_in_0_0_eta_V => tracks_in_0_0_eta_V,
                     tracks_in_0_1_eta_V => tracks_in_0_1_eta_V,
                     tracks_in_1_0_eta_V => tracks_in_1_0_eta_V,
                     tracks_in_1_1_eta_V => tracks_in_1_1_eta_V,
                     tracks_in_2_0_eta_V => tracks_in_2_0_eta_V,
                     tracks_in_2_1_eta_V => tracks_in_2_1_eta_V,
                     tracks_in_3_0_eta_V => tracks_in_3_0_eta_V,
                     tracks_in_3_1_eta_V => tracks_in_3_1_eta_V,
                     tracks_in_4_0_eta_V => tracks_in_4_0_eta_V,
                     tracks_in_4_1_eta_V => tracks_in_4_1_eta_V,
                     tracks_in_5_0_eta_V => tracks_in_5_0_eta_V,
                     tracks_in_5_1_eta_V => tracks_in_5_1_eta_V,
                     tracks_in_6_0_eta_V => tracks_in_6_0_eta_V,
                     tracks_in_6_1_eta_V => tracks_in_6_1_eta_V,
                     tracks_in_7_0_eta_V => tracks_in_7_0_eta_V,
                     tracks_in_7_1_eta_V => tracks_in_7_1_eta_V,
                     tracks_in_8_0_eta_V => tracks_in_8_0_eta_V,
                     tracks_in_8_1_eta_V => tracks_in_8_1_eta_V,
                     tracks_in_0_0_phi_V => tracks_in_0_0_phi_V,
                     tracks_in_0_1_phi_V => tracks_in_0_1_phi_V,
                     tracks_in_1_0_phi_V => tracks_in_1_0_phi_V,
                     tracks_in_1_1_phi_V => tracks_in_1_1_phi_V,
                     tracks_in_2_0_phi_V => tracks_in_2_0_phi_V,
                     tracks_in_2_1_phi_V => tracks_in_2_1_phi_V,
                     tracks_in_3_0_phi_V => tracks_in_3_0_phi_V,
                     tracks_in_3_1_phi_V => tracks_in_3_1_phi_V,
                     tracks_in_4_0_phi_V => tracks_in_4_0_phi_V,
                     tracks_in_4_1_phi_V => tracks_in_4_1_phi_V,
                     tracks_in_5_0_phi_V => tracks_in_5_0_phi_V,
                     tracks_in_5_1_phi_V => tracks_in_5_1_phi_V,
                     tracks_in_6_0_phi_V => tracks_in_6_0_phi_V,
                     tracks_in_6_1_phi_V => tracks_in_6_1_phi_V,
                     tracks_in_7_0_phi_V => tracks_in_7_0_phi_V,
                     tracks_in_7_1_phi_V => tracks_in_7_1_phi_V,
                     tracks_in_8_0_phi_V => tracks_in_8_0_phi_V,
                     tracks_in_8_1_phi_V => tracks_in_8_1_phi_V,
                     tracks_in_0_0_rest_V => tracks_in_0_0_rest_V,
                     tracks_in_0_1_rest_V => tracks_in_0_1_rest_V,
                     tracks_in_1_0_rest_V => tracks_in_1_0_rest_V,
                     tracks_in_1_1_rest_V => tracks_in_1_1_rest_V,
                     tracks_in_2_0_rest_V => tracks_in_2_0_rest_V,
                     tracks_in_2_1_rest_V => tracks_in_2_1_rest_V,
                     tracks_in_3_0_rest_V => tracks_in_3_0_rest_V,
                     tracks_in_3_1_rest_V => tracks_in_3_1_rest_V,
                     tracks_in_4_0_rest_V => tracks_in_4_0_rest_V,
                     tracks_in_4_1_rest_V => tracks_in_4_1_rest_V,
                     tracks_in_5_0_rest_V => tracks_in_5_0_rest_V,
                     tracks_in_5_1_rest_V => tracks_in_5_1_rest_V,
                     tracks_in_6_0_rest_V => tracks_in_6_0_rest_V,
                     tracks_in_6_1_rest_V => tracks_in_6_1_rest_V,
                     tracks_in_7_0_rest_V => tracks_in_7_0_rest_V,
                     tracks_in_7_1_rest_V => tracks_in_7_1_rest_V,
                     tracks_in_8_0_rest_V => tracks_in_8_0_rest_V,
                     tracks_in_8_1_rest_V => tracks_in_8_1_rest_V,
                     fifo_in_0_0_pt_V => fifo_in(0*NFIFOS+0).pt,
                     fifo_in_0_1_pt_V => fifo_in(0*NFIFOS+1).pt,
                     fifo_in_0_2_pt_V => fifo_in(0*NFIFOS+2).pt,
                     fifo_in_0_3_pt_V => fifo_in(0*NFIFOS+3).pt,
                     fifo_in_0_4_pt_V => fifo_in(0*NFIFOS+4).pt,
                     fifo_in_0_5_pt_V => fifo_in(0*NFIFOS+5).pt,
                     fifo_in_0_0_eta_V => fifo_in(0*NFIFOS+0).eta,
                     fifo_in_0_1_eta_V => fifo_in(0*NFIFOS+1).eta,
                     fifo_in_0_2_eta_V => fifo_in(0*NFIFOS+2).eta,
                     fifo_in_0_3_eta_V => fifo_in(0*NFIFOS+3).eta,
                     fifo_in_0_4_eta_V => fifo_in(0*NFIFOS+4).eta,
                     fifo_in_0_5_eta_V => fifo_in(0*NFIFOS+5).eta,
                     fifo_in_0_0_phi_V => fifo_in(0*NFIFOS+0).phi,
                     fifo_in_0_1_phi_V => fifo_in(0*NFIFOS+1).phi,
                     fifo_in_0_2_phi_V => fifo_in(0*NFIFOS+2).phi,
                     fifo_in_0_3_phi_V => fifo_in(0*NFIFOS+3).phi,
                     fifo_in_0_4_phi_V => fifo_in(0*NFIFOS+4).phi,
                     fifo_in_0_5_phi_V => fifo_in(0*NFIFOS+5).phi,
                     fifo_in_0_0_rest_V => fifo_in(0*NFIFOS+0).rest,
                     fifo_in_0_1_rest_V => fifo_in(0*NFIFOS+1).rest,
                     fifo_in_0_2_rest_V => fifo_in(0*NFIFOS+2).rest,
                     fifo_in_0_3_rest_V => fifo_in(0*NFIFOS+3).rest,
                     fifo_in_0_4_rest_V => fifo_in(0*NFIFOS+4).rest,
                     fifo_in_0_5_rest_V => fifo_in(0*NFIFOS+5).rest,
                     fifo_in_1_0_pt_V => fifo_in(1*NFIFOS+0).pt,
                     fifo_in_1_1_pt_V => fifo_in(1*NFIFOS+1).pt,
                     fifo_in_1_2_pt_V => fifo_in(1*NFIFOS+2).pt,
                     fifo_in_1_3_pt_V => fifo_in(1*NFIFOS+3).pt,
                     fifo_in_1_4_pt_V => fifo_in(1*NFIFOS+4).pt,
                     fifo_in_1_5_pt_V => fifo_in(1*NFIFOS+5).pt,
                     fifo_in_1_0_eta_V => fifo_in(1*NFIFOS+0).eta,
                     fifo_in_1_1_eta_V => fifo_in(1*NFIFOS+1).eta,
                     fifo_in_1_2_eta_V => fifo_in(1*NFIFOS+2).eta,
                     fifo_in_1_3_eta_V => fifo_in(1*NFIFOS+3).eta,
                     fifo_in_1_4_eta_V => fifo_in(1*NFIFOS+4).eta,
                     fifo_in_1_5_eta_V => fifo_in(1*NFIFOS+5).eta,
                     fifo_in_1_0_phi_V => fifo_in(1*NFIFOS+0).phi,
                     fifo_in_1_1_phi_V => fifo_in(1*NFIFOS+1).phi,
                     fifo_in_1_2_phi_V => fifo_in(1*NFIFOS+2).phi,
                     fifo_in_1_3_phi_V => fifo_in(1*NFIFOS+3).phi,
                     fifo_in_1_4_phi_V => fifo_in(1*NFIFOS+4).phi,
                     fifo_in_1_5_phi_V => fifo_in(1*NFIFOS+5).phi,
                     fifo_in_1_0_rest_V => fifo_in(1*NFIFOS+0).rest,
                     fifo_in_1_1_rest_V => fifo_in(1*NFIFOS+1).rest,
                     fifo_in_1_2_rest_V => fifo_in(1*NFIFOS+2).rest,
                     fifo_in_1_3_rest_V => fifo_in(1*NFIFOS+3).rest,
                     fifo_in_1_4_rest_V => fifo_in(1*NFIFOS+4).rest,
                     fifo_in_1_5_rest_V => fifo_in(1*NFIFOS+5).rest,
                     fifo_in_2_0_pt_V => fifo_in(2*NFIFOS+0).pt,
                     fifo_in_2_1_pt_V => fifo_in(2*NFIFOS+1).pt,
                     fifo_in_2_2_pt_V => fifo_in(2*NFIFOS+2).pt,
                     fifo_in_2_3_pt_V => fifo_in(2*NFIFOS+3).pt,
                     fifo_in_2_4_pt_V => fifo_in(2*NFIFOS+4).pt,
                     fifo_in_2_5_pt_V => fifo_in(2*NFIFOS+5).pt,
                     fifo_in_2_0_eta_V => fifo_in(2*NFIFOS+0).eta,
                     fifo_in_2_1_eta_V => fifo_in(2*NFIFOS+1).eta,
                     fifo_in_2_2_eta_V => fifo_in(2*NFIFOS+2).eta,
                     fifo_in_2_3_eta_V => fifo_in(2*NFIFOS+3).eta,
                     fifo_in_2_4_eta_V => fifo_in(2*NFIFOS+4).eta,
                     fifo_in_2_5_eta_V => fifo_in(2*NFIFOS+5).eta,
                     fifo_in_2_0_phi_V => fifo_in(2*NFIFOS+0).phi,
                     fifo_in_2_1_phi_V => fifo_in(2*NFIFOS+1).phi,
                     fifo_in_2_2_phi_V => fifo_in(2*NFIFOS+2).phi,
                     fifo_in_2_3_phi_V => fifo_in(2*NFIFOS+3).phi,
                     fifo_in_2_4_phi_V => fifo_in(2*NFIFOS+4).phi,
                     fifo_in_2_5_phi_V => fifo_in(2*NFIFOS+5).phi,
                     fifo_in_2_0_rest_V => fifo_in(2*NFIFOS+0).rest,
                     fifo_in_2_1_rest_V => fifo_in(2*NFIFOS+1).rest,
                     fifo_in_2_2_rest_V => fifo_in(2*NFIFOS+2).rest,
                     fifo_in_2_3_rest_V => fifo_in(2*NFIFOS+3).rest,
                     fifo_in_2_4_rest_V => fifo_in(2*NFIFOS+4).rest,
                     fifo_in_2_5_rest_V => fifo_in(2*NFIFOS+5).rest,
                     fifo_in_3_0_pt_V => fifo_in(3*NFIFOS+0).pt,
                     fifo_in_3_1_pt_V => fifo_in(3*NFIFOS+1).pt,
                     fifo_in_3_2_pt_V => fifo_in(3*NFIFOS+2).pt,
                     fifo_in_3_3_pt_V => fifo_in(3*NFIFOS+3).pt,
                     fifo_in_3_4_pt_V => fifo_in(3*NFIFOS+4).pt,
                     fifo_in_3_5_pt_V => fifo_in(3*NFIFOS+5).pt,
                     fifo_in_3_0_eta_V => fifo_in(3*NFIFOS+0).eta,
                     fifo_in_3_1_eta_V => fifo_in(3*NFIFOS+1).eta,
                     fifo_in_3_2_eta_V => fifo_in(3*NFIFOS+2).eta,
                     fifo_in_3_3_eta_V => fifo_in(3*NFIFOS+3).eta,
                     fifo_in_3_4_eta_V => fifo_in(3*NFIFOS+4).eta,
                     fifo_in_3_5_eta_V => fifo_in(3*NFIFOS+5).eta,
                     fifo_in_3_0_phi_V => fifo_in(3*NFIFOS+0).phi,
                     fifo_in_3_1_phi_V => fifo_in(3*NFIFOS+1).phi,
                     fifo_in_3_2_phi_V => fifo_in(3*NFIFOS+2).phi,
                     fifo_in_3_3_phi_V => fifo_in(3*NFIFOS+3).phi,
                     fifo_in_3_4_phi_V => fifo_in(3*NFIFOS+4).phi,
                     fifo_in_3_5_phi_V => fifo_in(3*NFIFOS+5).phi,
                     fifo_in_3_0_rest_V => fifo_in(3*NFIFOS+0).rest,
                     fifo_in_3_1_rest_V => fifo_in(3*NFIFOS+1).rest,
                     fifo_in_3_2_rest_V => fifo_in(3*NFIFOS+2).rest,
                     fifo_in_3_3_rest_V => fifo_in(3*NFIFOS+3).rest,
                     fifo_in_3_4_rest_V => fifo_in(3*NFIFOS+4).rest,
                     fifo_in_3_5_rest_V => fifo_in(3*NFIFOS+5).rest,
                     fifo_in_4_0_pt_V => fifo_in(4*NFIFOS+0).pt,
                     fifo_in_4_1_pt_V => fifo_in(4*NFIFOS+1).pt,
                     fifo_in_4_2_pt_V => fifo_in(4*NFIFOS+2).pt,
                     fifo_in_4_3_pt_V => fifo_in(4*NFIFOS+3).pt,
                     fifo_in_4_4_pt_V => fifo_in(4*NFIFOS+4).pt,
                     fifo_in_4_5_pt_V => fifo_in(4*NFIFOS+5).pt,
                     fifo_in_4_0_eta_V => fifo_in(4*NFIFOS+0).eta,
                     fifo_in_4_1_eta_V => fifo_in(4*NFIFOS+1).eta,
                     fifo_in_4_2_eta_V => fifo_in(4*NFIFOS+2).eta,
                     fifo_in_4_3_eta_V => fifo_in(4*NFIFOS+3).eta,
                     fifo_in_4_4_eta_V => fifo_in(4*NFIFOS+4).eta,
                     fifo_in_4_5_eta_V => fifo_in(4*NFIFOS+5).eta,
                     fifo_in_4_0_phi_V => fifo_in(4*NFIFOS+0).phi,
                     fifo_in_4_1_phi_V => fifo_in(4*NFIFOS+1).phi,
                     fifo_in_4_2_phi_V => fifo_in(4*NFIFOS+2).phi,
                     fifo_in_4_3_phi_V => fifo_in(4*NFIFOS+3).phi,
                     fifo_in_4_4_phi_V => fifo_in(4*NFIFOS+4).phi,
                     fifo_in_4_5_phi_V => fifo_in(4*NFIFOS+5).phi,
                     fifo_in_4_0_rest_V => fifo_in(4*NFIFOS+0).rest,
                     fifo_in_4_1_rest_V => fifo_in(4*NFIFOS+1).rest,
                     fifo_in_4_2_rest_V => fifo_in(4*NFIFOS+2).rest,
                     fifo_in_4_3_rest_V => fifo_in(4*NFIFOS+3).rest,
                     fifo_in_4_4_rest_V => fifo_in(4*NFIFOS+4).rest,
                     fifo_in_4_5_rest_V => fifo_in(4*NFIFOS+5).rest,
                     fifo_in_5_0_pt_V => fifo_in(5*NFIFOS+0).pt,
                     fifo_in_5_1_pt_V => fifo_in(5*NFIFOS+1).pt,
                     fifo_in_5_2_pt_V => fifo_in(5*NFIFOS+2).pt,
                     fifo_in_5_3_pt_V => fifo_in(5*NFIFOS+3).pt,
                     fifo_in_5_4_pt_V => fifo_in(5*NFIFOS+4).pt,
                     fifo_in_5_5_pt_V => fifo_in(5*NFIFOS+5).pt,
                     fifo_in_5_0_eta_V => fifo_in(5*NFIFOS+0).eta,
                     fifo_in_5_1_eta_V => fifo_in(5*NFIFOS+1).eta,
                     fifo_in_5_2_eta_V => fifo_in(5*NFIFOS+2).eta,
                     fifo_in_5_3_eta_V => fifo_in(5*NFIFOS+3).eta,
                     fifo_in_5_4_eta_V => fifo_in(5*NFIFOS+4).eta,
                     fifo_in_5_5_eta_V => fifo_in(5*NFIFOS+5).eta,
                     fifo_in_5_0_phi_V => fifo_in(5*NFIFOS+0).phi,
                     fifo_in_5_1_phi_V => fifo_in(5*NFIFOS+1).phi,
                     fifo_in_5_2_phi_V => fifo_in(5*NFIFOS+2).phi,
                     fifo_in_5_3_phi_V => fifo_in(5*NFIFOS+3).phi,
                     fifo_in_5_4_phi_V => fifo_in(5*NFIFOS+4).phi,
                     fifo_in_5_5_phi_V => fifo_in(5*NFIFOS+5).phi,
                     fifo_in_5_0_rest_V => fifo_in(5*NFIFOS+0).rest,
                     fifo_in_5_1_rest_V => fifo_in(5*NFIFOS+1).rest,
                     fifo_in_5_2_rest_V => fifo_in(5*NFIFOS+2).rest,
                     fifo_in_5_3_rest_V => fifo_in(5*NFIFOS+3).rest,
                     fifo_in_5_4_rest_V => fifo_in(5*NFIFOS+4).rest,
                     fifo_in_5_5_rest_V => fifo_in(5*NFIFOS+5).rest,
                     fifo_in_6_0_pt_V => fifo_in(6*NFIFOS+0).pt,
                     fifo_in_6_1_pt_V => fifo_in(6*NFIFOS+1).pt,
                     fifo_in_6_2_pt_V => fifo_in(6*NFIFOS+2).pt,
                     fifo_in_6_3_pt_V => fifo_in(6*NFIFOS+3).pt,
                     fifo_in_6_4_pt_V => fifo_in(6*NFIFOS+4).pt,
                     fifo_in_6_5_pt_V => fifo_in(6*NFIFOS+5).pt,
                     fifo_in_6_0_eta_V => fifo_in(6*NFIFOS+0).eta,
                     fifo_in_6_1_eta_V => fifo_in(6*NFIFOS+1).eta,
                     fifo_in_6_2_eta_V => fifo_in(6*NFIFOS+2).eta,
                     fifo_in_6_3_eta_V => fifo_in(6*NFIFOS+3).eta,
                     fifo_in_6_4_eta_V => fifo_in(6*NFIFOS+4).eta,
                     fifo_in_6_5_eta_V => fifo_in(6*NFIFOS+5).eta,
                     fifo_in_6_0_phi_V => fifo_in(6*NFIFOS+0).phi,
                     fifo_in_6_1_phi_V => fifo_in(6*NFIFOS+1).phi,
                     fifo_in_6_2_phi_V => fifo_in(6*NFIFOS+2).phi,
                     fifo_in_6_3_phi_V => fifo_in(6*NFIFOS+3).phi,
                     fifo_in_6_4_phi_V => fifo_in(6*NFIFOS+4).phi,
                     fifo_in_6_5_phi_V => fifo_in(6*NFIFOS+5).phi,
                     fifo_in_6_0_rest_V => fifo_in(6*NFIFOS+0).rest,
                     fifo_in_6_1_rest_V => fifo_in(6*NFIFOS+1).rest,
                     fifo_in_6_2_rest_V => fifo_in(6*NFIFOS+2).rest,
                     fifo_in_6_3_rest_V => fifo_in(6*NFIFOS+3).rest,
                     fifo_in_6_4_rest_V => fifo_in(6*NFIFOS+4).rest,
                     fifo_in_6_5_rest_V => fifo_in(6*NFIFOS+5).rest,
                     fifo_in_7_0_pt_V => fifo_in(7*NFIFOS+0).pt,
                     fifo_in_7_1_pt_V => fifo_in(7*NFIFOS+1).pt,
                     fifo_in_7_2_pt_V => fifo_in(7*NFIFOS+2).pt,
                     fifo_in_7_3_pt_V => fifo_in(7*NFIFOS+3).pt,
                     fifo_in_7_4_pt_V => fifo_in(7*NFIFOS+4).pt,
                     fifo_in_7_5_pt_V => fifo_in(7*NFIFOS+5).pt,
                     fifo_in_7_0_eta_V => fifo_in(7*NFIFOS+0).eta,
                     fifo_in_7_1_eta_V => fifo_in(7*NFIFOS+1).eta,
                     fifo_in_7_2_eta_V => fifo_in(7*NFIFOS+2).eta,
                     fifo_in_7_3_eta_V => fifo_in(7*NFIFOS+3).eta,
                     fifo_in_7_4_eta_V => fifo_in(7*NFIFOS+4).eta,
                     fifo_in_7_5_eta_V => fifo_in(7*NFIFOS+5).eta,
                     fifo_in_7_0_phi_V => fifo_in(7*NFIFOS+0).phi,
                     fifo_in_7_1_phi_V => fifo_in(7*NFIFOS+1).phi,
                     fifo_in_7_2_phi_V => fifo_in(7*NFIFOS+2).phi,
                     fifo_in_7_3_phi_V => fifo_in(7*NFIFOS+3).phi,
                     fifo_in_7_4_phi_V => fifo_in(7*NFIFOS+4).phi,
                     fifo_in_7_5_phi_V => fifo_in(7*NFIFOS+5).phi,
                     fifo_in_7_0_rest_V => fifo_in(7*NFIFOS+0).rest,
                     fifo_in_7_1_rest_V => fifo_in(7*NFIFOS+1).rest,
                     fifo_in_7_2_rest_V => fifo_in(7*NFIFOS+2).rest,
                     fifo_in_7_3_rest_V => fifo_in(7*NFIFOS+3).rest,
                     fifo_in_7_4_rest_V => fifo_in(7*NFIFOS+4).rest,
                     fifo_in_7_5_rest_V => fifo_in(7*NFIFOS+5).rest,
                     fifo_in_8_0_pt_V => fifo_in(8*NFIFOS+0).pt,
                     fifo_in_8_1_pt_V => fifo_in(8*NFIFOS+1).pt,
                     fifo_in_8_2_pt_V => fifo_in(8*NFIFOS+2).pt,
                     fifo_in_8_3_pt_V => fifo_in(8*NFIFOS+3).pt,
                     fifo_in_8_4_pt_V => fifo_in(8*NFIFOS+4).pt,
                     fifo_in_8_5_pt_V => fifo_in(8*NFIFOS+5).pt,
                     fifo_in_8_0_eta_V => fifo_in(8*NFIFOS+0).eta,
                     fifo_in_8_1_eta_V => fifo_in(8*NFIFOS+1).eta,
                     fifo_in_8_2_eta_V => fifo_in(8*NFIFOS+2).eta,
                     fifo_in_8_3_eta_V => fifo_in(8*NFIFOS+3).eta,
                     fifo_in_8_4_eta_V => fifo_in(8*NFIFOS+4).eta,
                     fifo_in_8_5_eta_V => fifo_in(8*NFIFOS+5).eta,
                     fifo_in_8_0_phi_V => fifo_in(8*NFIFOS+0).phi,
                     fifo_in_8_1_phi_V => fifo_in(8*NFIFOS+1).phi,
                     fifo_in_8_2_phi_V => fifo_in(8*NFIFOS+2).phi,
                     fifo_in_8_3_phi_V => fifo_in(8*NFIFOS+3).phi,
                     fifo_in_8_4_phi_V => fifo_in(8*NFIFOS+4).phi,
                     fifo_in_8_5_phi_V => fifo_in(8*NFIFOS+5).phi,
                     fifo_in_8_0_rest_V => fifo_in(8*NFIFOS+0).rest,
                     fifo_in_8_1_rest_V => fifo_in(8*NFIFOS+1).rest,
                     fifo_in_8_2_rest_V => fifo_in(8*NFIFOS+2).rest,
                     fifo_in_8_3_rest_V => fifo_in(8*NFIFOS+3).rest,
                     fifo_in_8_4_rest_V => fifo_in(8*NFIFOS+4).rest,
                     fifo_in_8_5_rest_V => fifo_in(8*NFIFOS+5).rest,
                     fifo_write_0_0 => fifo_in_write(0*NFIFOS+0),
                     fifo_write_0_1 => fifo_in_write(0*NFIFOS+1),
                     fifo_write_0_2 => fifo_in_write(0*NFIFOS+2),
                     fifo_write_0_3 => fifo_in_write(0*NFIFOS+3),
                     fifo_write_0_4 => fifo_in_write(0*NFIFOS+4),
                     fifo_write_0_5 => fifo_in_write(0*NFIFOS+5),
                     fifo_write_1_0 => fifo_in_write(1*NFIFOS+0),
                     fifo_write_1_1 => fifo_in_write(1*NFIFOS+1),
                     fifo_write_1_2 => fifo_in_write(1*NFIFOS+2),
                     fifo_write_1_3 => fifo_in_write(1*NFIFOS+3),
                     fifo_write_1_4 => fifo_in_write(1*NFIFOS+4),
                     fifo_write_1_5 => fifo_in_write(1*NFIFOS+5),
                     fifo_write_2_0 => fifo_in_write(2*NFIFOS+0),
                     fifo_write_2_1 => fifo_in_write(2*NFIFOS+1),
                     fifo_write_2_2 => fifo_in_write(2*NFIFOS+2),
                     fifo_write_2_3 => fifo_in_write(2*NFIFOS+3),
                     fifo_write_2_4 => fifo_in_write(2*NFIFOS+4),
                     fifo_write_2_5 => fifo_in_write(2*NFIFOS+5),
                     fifo_write_3_0 => fifo_in_write(3*NFIFOS+0),
                     fifo_write_3_1 => fifo_in_write(3*NFIFOS+1),
                     fifo_write_3_2 => fifo_in_write(3*NFIFOS+2),
                     fifo_write_3_3 => fifo_in_write(3*NFIFOS+3),
                     fifo_write_3_4 => fifo_in_write(3*NFIFOS+4),
                     fifo_write_3_5 => fifo_in_write(3*NFIFOS+5),
                     fifo_write_4_0 => fifo_in_write(4*NFIFOS+0),
                     fifo_write_4_1 => fifo_in_write(4*NFIFOS+1),
                     fifo_write_4_2 => fifo_in_write(4*NFIFOS+2),
                     fifo_write_4_3 => fifo_in_write(4*NFIFOS+3),
                     fifo_write_4_4 => fifo_in_write(4*NFIFOS+4),
                     fifo_write_4_5 => fifo_in_write(4*NFIFOS+5),
                     fifo_write_5_0 => fifo_in_write(5*NFIFOS+0),
                     fifo_write_5_1 => fifo_in_write(5*NFIFOS+1),
                     fifo_write_5_2 => fifo_in_write(5*NFIFOS+2),
                     fifo_write_5_3 => fifo_in_write(5*NFIFOS+3),
                     fifo_write_5_4 => fifo_in_write(5*NFIFOS+4),
                     fifo_write_5_5 => fifo_in_write(5*NFIFOS+5),
                     fifo_write_6_0 => fifo_in_write(6*NFIFOS+0),
                     fifo_write_6_1 => fifo_in_write(6*NFIFOS+1),
                     fifo_write_6_2 => fifo_in_write(6*NFIFOS+2),
                     fifo_write_6_3 => fifo_in_write(6*NFIFOS+3),
                     fifo_write_6_4 => fifo_in_write(6*NFIFOS+4),
                     fifo_write_6_5 => fifo_in_write(6*NFIFOS+5),
                     fifo_write_7_0 => fifo_in_write(7*NFIFOS+0),
                     fifo_write_7_1 => fifo_in_write(7*NFIFOS+1),
                     fifo_write_7_2 => fifo_in_write(7*NFIFOS+2),
                     fifo_write_7_3 => fifo_in_write(7*NFIFOS+3),
                     fifo_write_7_4 => fifo_in_write(7*NFIFOS+4),
                     fifo_write_7_5 => fifo_in_write(7*NFIFOS+5),
                     fifo_write_8_0 => fifo_in_write(8*NFIFOS+0),
                     fifo_write_8_1 => fifo_in_write(8*NFIFOS+1),
                     fifo_write_8_2 => fifo_in_write(8*NFIFOS+2),
                     fifo_write_8_3 => fifo_in_write(8*NFIFOS+3),
                     fifo_write_8_4 => fifo_in_write(8*NFIFOS+4),
                     fifo_write_8_5 => fifo_in_write(8*NFIFOS+5)
                    );

    fifo_slice : entity work.router_fifo_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     newevent => newevent_del,
                     fifo_in_0_0_pt_V => fifo_in(0*NFIFOS+0).pt,
                     fifo_in_0_1_pt_V => fifo_in(0*NFIFOS+1).pt,
                     fifo_in_0_2_pt_V => fifo_in(0*NFIFOS+2).pt,
                     fifo_in_0_3_pt_V => fifo_in(0*NFIFOS+3).pt,
                     fifo_in_0_4_pt_V => fifo_in(0*NFIFOS+4).pt,
                     fifo_in_0_5_pt_V => fifo_in(0*NFIFOS+5).pt,
                     fifo_in_0_0_eta_V => fifo_in(0*NFIFOS+0).eta,
                     fifo_in_0_1_eta_V => fifo_in(0*NFIFOS+1).eta,
                     fifo_in_0_2_eta_V => fifo_in(0*NFIFOS+2).eta,
                     fifo_in_0_3_eta_V => fifo_in(0*NFIFOS+3).eta,
                     fifo_in_0_4_eta_V => fifo_in(0*NFIFOS+4).eta,
                     fifo_in_0_5_eta_V => fifo_in(0*NFIFOS+5).eta,
                     fifo_in_0_0_phi_V => fifo_in(0*NFIFOS+0).phi,
                     fifo_in_0_1_phi_V => fifo_in(0*NFIFOS+1).phi,
                     fifo_in_0_2_phi_V => fifo_in(0*NFIFOS+2).phi,
                     fifo_in_0_3_phi_V => fifo_in(0*NFIFOS+3).phi,
                     fifo_in_0_4_phi_V => fifo_in(0*NFIFOS+4).phi,
                     fifo_in_0_5_phi_V => fifo_in(0*NFIFOS+5).phi,
                     fifo_in_0_0_rest_V => fifo_in(0*NFIFOS+0).rest,
                     fifo_in_0_1_rest_V => fifo_in(0*NFIFOS+1).rest,
                     fifo_in_0_2_rest_V => fifo_in(0*NFIFOS+2).rest,
                     fifo_in_0_3_rest_V => fifo_in(0*NFIFOS+3).rest,
                     fifo_in_0_4_rest_V => fifo_in(0*NFIFOS+4).rest,
                     fifo_in_0_5_rest_V => fifo_in(0*NFIFOS+5).rest,
                     fifo_in_1_0_pt_V => fifo_in(1*NFIFOS+0).pt,
                     fifo_in_1_1_pt_V => fifo_in(1*NFIFOS+1).pt,
                     fifo_in_1_2_pt_V => fifo_in(1*NFIFOS+2).pt,
                     fifo_in_1_3_pt_V => fifo_in(1*NFIFOS+3).pt,
                     fifo_in_1_4_pt_V => fifo_in(1*NFIFOS+4).pt,
                     fifo_in_1_5_pt_V => fifo_in(1*NFIFOS+5).pt,
                     fifo_in_1_0_eta_V => fifo_in(1*NFIFOS+0).eta,
                     fifo_in_1_1_eta_V => fifo_in(1*NFIFOS+1).eta,
                     fifo_in_1_2_eta_V => fifo_in(1*NFIFOS+2).eta,
                     fifo_in_1_3_eta_V => fifo_in(1*NFIFOS+3).eta,
                     fifo_in_1_4_eta_V => fifo_in(1*NFIFOS+4).eta,
                     fifo_in_1_5_eta_V => fifo_in(1*NFIFOS+5).eta,
                     fifo_in_1_0_phi_V => fifo_in(1*NFIFOS+0).phi,
                     fifo_in_1_1_phi_V => fifo_in(1*NFIFOS+1).phi,
                     fifo_in_1_2_phi_V => fifo_in(1*NFIFOS+2).phi,
                     fifo_in_1_3_phi_V => fifo_in(1*NFIFOS+3).phi,
                     fifo_in_1_4_phi_V => fifo_in(1*NFIFOS+4).phi,
                     fifo_in_1_5_phi_V => fifo_in(1*NFIFOS+5).phi,
                     fifo_in_1_0_rest_V => fifo_in(1*NFIFOS+0).rest,
                     fifo_in_1_1_rest_V => fifo_in(1*NFIFOS+1).rest,
                     fifo_in_1_2_rest_V => fifo_in(1*NFIFOS+2).rest,
                     fifo_in_1_3_rest_V => fifo_in(1*NFIFOS+3).rest,
                     fifo_in_1_4_rest_V => fifo_in(1*NFIFOS+4).rest,
                     fifo_in_1_5_rest_V => fifo_in(1*NFIFOS+5).rest,
                     fifo_in_2_0_pt_V => fifo_in(2*NFIFOS+0).pt,
                     fifo_in_2_1_pt_V => fifo_in(2*NFIFOS+1).pt,
                     fifo_in_2_2_pt_V => fifo_in(2*NFIFOS+2).pt,
                     fifo_in_2_3_pt_V => fifo_in(2*NFIFOS+3).pt,
                     fifo_in_2_4_pt_V => fifo_in(2*NFIFOS+4).pt,
                     fifo_in_2_5_pt_V => fifo_in(2*NFIFOS+5).pt,
                     fifo_in_2_0_eta_V => fifo_in(2*NFIFOS+0).eta,
                     fifo_in_2_1_eta_V => fifo_in(2*NFIFOS+1).eta,
                     fifo_in_2_2_eta_V => fifo_in(2*NFIFOS+2).eta,
                     fifo_in_2_3_eta_V => fifo_in(2*NFIFOS+3).eta,
                     fifo_in_2_4_eta_V => fifo_in(2*NFIFOS+4).eta,
                     fifo_in_2_5_eta_V => fifo_in(2*NFIFOS+5).eta,
                     fifo_in_2_0_phi_V => fifo_in(2*NFIFOS+0).phi,
                     fifo_in_2_1_phi_V => fifo_in(2*NFIFOS+1).phi,
                     fifo_in_2_2_phi_V => fifo_in(2*NFIFOS+2).phi,
                     fifo_in_2_3_phi_V => fifo_in(2*NFIFOS+3).phi,
                     fifo_in_2_4_phi_V => fifo_in(2*NFIFOS+4).phi,
                     fifo_in_2_5_phi_V => fifo_in(2*NFIFOS+5).phi,
                     fifo_in_2_0_rest_V => fifo_in(2*NFIFOS+0).rest,
                     fifo_in_2_1_rest_V => fifo_in(2*NFIFOS+1).rest,
                     fifo_in_2_2_rest_V => fifo_in(2*NFIFOS+2).rest,
                     fifo_in_2_3_rest_V => fifo_in(2*NFIFOS+3).rest,
                     fifo_in_2_4_rest_V => fifo_in(2*NFIFOS+4).rest,
                     fifo_in_2_5_rest_V => fifo_in(2*NFIFOS+5).rest,
                     fifo_in_3_0_pt_V => fifo_in(3*NFIFOS+0).pt,
                     fifo_in_3_1_pt_V => fifo_in(3*NFIFOS+1).pt,
                     fifo_in_3_2_pt_V => fifo_in(3*NFIFOS+2).pt,
                     fifo_in_3_3_pt_V => fifo_in(3*NFIFOS+3).pt,
                     fifo_in_3_4_pt_V => fifo_in(3*NFIFOS+4).pt,
                     fifo_in_3_5_pt_V => fifo_in(3*NFIFOS+5).pt,
                     fifo_in_3_0_eta_V => fifo_in(3*NFIFOS+0).eta,
                     fifo_in_3_1_eta_V => fifo_in(3*NFIFOS+1).eta,
                     fifo_in_3_2_eta_V => fifo_in(3*NFIFOS+2).eta,
                     fifo_in_3_3_eta_V => fifo_in(3*NFIFOS+3).eta,
                     fifo_in_3_4_eta_V => fifo_in(3*NFIFOS+4).eta,
                     fifo_in_3_5_eta_V => fifo_in(3*NFIFOS+5).eta,
                     fifo_in_3_0_phi_V => fifo_in(3*NFIFOS+0).phi,
                     fifo_in_3_1_phi_V => fifo_in(3*NFIFOS+1).phi,
                     fifo_in_3_2_phi_V => fifo_in(3*NFIFOS+2).phi,
                     fifo_in_3_3_phi_V => fifo_in(3*NFIFOS+3).phi,
                     fifo_in_3_4_phi_V => fifo_in(3*NFIFOS+4).phi,
                     fifo_in_3_5_phi_V => fifo_in(3*NFIFOS+5).phi,
                     fifo_in_3_0_rest_V => fifo_in(3*NFIFOS+0).rest,
                     fifo_in_3_1_rest_V => fifo_in(3*NFIFOS+1).rest,
                     fifo_in_3_2_rest_V => fifo_in(3*NFIFOS+2).rest,
                     fifo_in_3_3_rest_V => fifo_in(3*NFIFOS+3).rest,
                     fifo_in_3_4_rest_V => fifo_in(3*NFIFOS+4).rest,
                     fifo_in_3_5_rest_V => fifo_in(3*NFIFOS+5).rest,
                     fifo_in_4_0_pt_V => fifo_in(4*NFIFOS+0).pt,
                     fifo_in_4_1_pt_V => fifo_in(4*NFIFOS+1).pt,
                     fifo_in_4_2_pt_V => fifo_in(4*NFIFOS+2).pt,
                     fifo_in_4_3_pt_V => fifo_in(4*NFIFOS+3).pt,
                     fifo_in_4_4_pt_V => fifo_in(4*NFIFOS+4).pt,
                     fifo_in_4_5_pt_V => fifo_in(4*NFIFOS+5).pt,
                     fifo_in_4_0_eta_V => fifo_in(4*NFIFOS+0).eta,
                     fifo_in_4_1_eta_V => fifo_in(4*NFIFOS+1).eta,
                     fifo_in_4_2_eta_V => fifo_in(4*NFIFOS+2).eta,
                     fifo_in_4_3_eta_V => fifo_in(4*NFIFOS+3).eta,
                     fifo_in_4_4_eta_V => fifo_in(4*NFIFOS+4).eta,
                     fifo_in_4_5_eta_V => fifo_in(4*NFIFOS+5).eta,
                     fifo_in_4_0_phi_V => fifo_in(4*NFIFOS+0).phi,
                     fifo_in_4_1_phi_V => fifo_in(4*NFIFOS+1).phi,
                     fifo_in_4_2_phi_V => fifo_in(4*NFIFOS+2).phi,
                     fifo_in_4_3_phi_V => fifo_in(4*NFIFOS+3).phi,
                     fifo_in_4_4_phi_V => fifo_in(4*NFIFOS+4).phi,
                     fifo_in_4_5_phi_V => fifo_in(4*NFIFOS+5).phi,
                     fifo_in_4_0_rest_V => fifo_in(4*NFIFOS+0).rest,
                     fifo_in_4_1_rest_V => fifo_in(4*NFIFOS+1).rest,
                     fifo_in_4_2_rest_V => fifo_in(4*NFIFOS+2).rest,
                     fifo_in_4_3_rest_V => fifo_in(4*NFIFOS+3).rest,
                     fifo_in_4_4_rest_V => fifo_in(4*NFIFOS+4).rest,
                     fifo_in_4_5_rest_V => fifo_in(4*NFIFOS+5).rest,
                     fifo_in_5_0_pt_V => fifo_in(5*NFIFOS+0).pt,
                     fifo_in_5_1_pt_V => fifo_in(5*NFIFOS+1).pt,
                     fifo_in_5_2_pt_V => fifo_in(5*NFIFOS+2).pt,
                     fifo_in_5_3_pt_V => fifo_in(5*NFIFOS+3).pt,
                     fifo_in_5_4_pt_V => fifo_in(5*NFIFOS+4).pt,
                     fifo_in_5_5_pt_V => fifo_in(5*NFIFOS+5).pt,
                     fifo_in_5_0_eta_V => fifo_in(5*NFIFOS+0).eta,
                     fifo_in_5_1_eta_V => fifo_in(5*NFIFOS+1).eta,
                     fifo_in_5_2_eta_V => fifo_in(5*NFIFOS+2).eta,
                     fifo_in_5_3_eta_V => fifo_in(5*NFIFOS+3).eta,
                     fifo_in_5_4_eta_V => fifo_in(5*NFIFOS+4).eta,
                     fifo_in_5_5_eta_V => fifo_in(5*NFIFOS+5).eta,
                     fifo_in_5_0_phi_V => fifo_in(5*NFIFOS+0).phi,
                     fifo_in_5_1_phi_V => fifo_in(5*NFIFOS+1).phi,
                     fifo_in_5_2_phi_V => fifo_in(5*NFIFOS+2).phi,
                     fifo_in_5_3_phi_V => fifo_in(5*NFIFOS+3).phi,
                     fifo_in_5_4_phi_V => fifo_in(5*NFIFOS+4).phi,
                     fifo_in_5_5_phi_V => fifo_in(5*NFIFOS+5).phi,
                     fifo_in_5_0_rest_V => fifo_in(5*NFIFOS+0).rest,
                     fifo_in_5_1_rest_V => fifo_in(5*NFIFOS+1).rest,
                     fifo_in_5_2_rest_V => fifo_in(5*NFIFOS+2).rest,
                     fifo_in_5_3_rest_V => fifo_in(5*NFIFOS+3).rest,
                     fifo_in_5_4_rest_V => fifo_in(5*NFIFOS+4).rest,
                     fifo_in_5_5_rest_V => fifo_in(5*NFIFOS+5).rest,
                     fifo_in_6_0_pt_V => fifo_in(6*NFIFOS+0).pt,
                     fifo_in_6_1_pt_V => fifo_in(6*NFIFOS+1).pt,
                     fifo_in_6_2_pt_V => fifo_in(6*NFIFOS+2).pt,
                     fifo_in_6_3_pt_V => fifo_in(6*NFIFOS+3).pt,
                     fifo_in_6_4_pt_V => fifo_in(6*NFIFOS+4).pt,
                     fifo_in_6_5_pt_V => fifo_in(6*NFIFOS+5).pt,
                     fifo_in_6_0_eta_V => fifo_in(6*NFIFOS+0).eta,
                     fifo_in_6_1_eta_V => fifo_in(6*NFIFOS+1).eta,
                     fifo_in_6_2_eta_V => fifo_in(6*NFIFOS+2).eta,
                     fifo_in_6_3_eta_V => fifo_in(6*NFIFOS+3).eta,
                     fifo_in_6_4_eta_V => fifo_in(6*NFIFOS+4).eta,
                     fifo_in_6_5_eta_V => fifo_in(6*NFIFOS+5).eta,
                     fifo_in_6_0_phi_V => fifo_in(6*NFIFOS+0).phi,
                     fifo_in_6_1_phi_V => fifo_in(6*NFIFOS+1).phi,
                     fifo_in_6_2_phi_V => fifo_in(6*NFIFOS+2).phi,
                     fifo_in_6_3_phi_V => fifo_in(6*NFIFOS+3).phi,
                     fifo_in_6_4_phi_V => fifo_in(6*NFIFOS+4).phi,
                     fifo_in_6_5_phi_V => fifo_in(6*NFIFOS+5).phi,
                     fifo_in_6_0_rest_V => fifo_in(6*NFIFOS+0).rest,
                     fifo_in_6_1_rest_V => fifo_in(6*NFIFOS+1).rest,
                     fifo_in_6_2_rest_V => fifo_in(6*NFIFOS+2).rest,
                     fifo_in_6_3_rest_V => fifo_in(6*NFIFOS+3).rest,
                     fifo_in_6_4_rest_V => fifo_in(6*NFIFOS+4).rest,
                     fifo_in_6_5_rest_V => fifo_in(6*NFIFOS+5).rest,
                     fifo_in_7_0_pt_V => fifo_in(7*NFIFOS+0).pt,
                     fifo_in_7_1_pt_V => fifo_in(7*NFIFOS+1).pt,
                     fifo_in_7_2_pt_V => fifo_in(7*NFIFOS+2).pt,
                     fifo_in_7_3_pt_V => fifo_in(7*NFIFOS+3).pt,
                     fifo_in_7_4_pt_V => fifo_in(7*NFIFOS+4).pt,
                     fifo_in_7_5_pt_V => fifo_in(7*NFIFOS+5).pt,
                     fifo_in_7_0_eta_V => fifo_in(7*NFIFOS+0).eta,
                     fifo_in_7_1_eta_V => fifo_in(7*NFIFOS+1).eta,
                     fifo_in_7_2_eta_V => fifo_in(7*NFIFOS+2).eta,
                     fifo_in_7_3_eta_V => fifo_in(7*NFIFOS+3).eta,
                     fifo_in_7_4_eta_V => fifo_in(7*NFIFOS+4).eta,
                     fifo_in_7_5_eta_V => fifo_in(7*NFIFOS+5).eta,
                     fifo_in_7_0_phi_V => fifo_in(7*NFIFOS+0).phi,
                     fifo_in_7_1_phi_V => fifo_in(7*NFIFOS+1).phi,
                     fifo_in_7_2_phi_V => fifo_in(7*NFIFOS+2).phi,
                     fifo_in_7_3_phi_V => fifo_in(7*NFIFOS+3).phi,
                     fifo_in_7_4_phi_V => fifo_in(7*NFIFOS+4).phi,
                     fifo_in_7_5_phi_V => fifo_in(7*NFIFOS+5).phi,
                     fifo_in_7_0_rest_V => fifo_in(7*NFIFOS+0).rest,
                     fifo_in_7_1_rest_V => fifo_in(7*NFIFOS+1).rest,
                     fifo_in_7_2_rest_V => fifo_in(7*NFIFOS+2).rest,
                     fifo_in_7_3_rest_V => fifo_in(7*NFIFOS+3).rest,
                     fifo_in_7_4_rest_V => fifo_in(7*NFIFOS+4).rest,
                     fifo_in_7_5_rest_V => fifo_in(7*NFIFOS+5).rest,
                     fifo_in_8_0_pt_V => fifo_in(8*NFIFOS+0).pt,
                     fifo_in_8_1_pt_V => fifo_in(8*NFIFOS+1).pt,
                     fifo_in_8_2_pt_V => fifo_in(8*NFIFOS+2).pt,
                     fifo_in_8_3_pt_V => fifo_in(8*NFIFOS+3).pt,
                     fifo_in_8_4_pt_V => fifo_in(8*NFIFOS+4).pt,
                     fifo_in_8_5_pt_V => fifo_in(8*NFIFOS+5).pt,
                     fifo_in_8_0_eta_V => fifo_in(8*NFIFOS+0).eta,
                     fifo_in_8_1_eta_V => fifo_in(8*NFIFOS+1).eta,
                     fifo_in_8_2_eta_V => fifo_in(8*NFIFOS+2).eta,
                     fifo_in_8_3_eta_V => fifo_in(8*NFIFOS+3).eta,
                     fifo_in_8_4_eta_V => fifo_in(8*NFIFOS+4).eta,
                     fifo_in_8_5_eta_V => fifo_in(8*NFIFOS+5).eta,
                     fifo_in_8_0_phi_V => fifo_in(8*NFIFOS+0).phi,
                     fifo_in_8_1_phi_V => fifo_in(8*NFIFOS+1).phi,
                     fifo_in_8_2_phi_V => fifo_in(8*NFIFOS+2).phi,
                     fifo_in_8_3_phi_V => fifo_in(8*NFIFOS+3).phi,
                     fifo_in_8_4_phi_V => fifo_in(8*NFIFOS+4).phi,
                     fifo_in_8_5_phi_V => fifo_in(8*NFIFOS+5).phi,
                     fifo_in_8_0_rest_V => fifo_in(8*NFIFOS+0).rest,
                     fifo_in_8_1_rest_V => fifo_in(8*NFIFOS+1).rest,
                     fifo_in_8_2_rest_V => fifo_in(8*NFIFOS+2).rest,
                     fifo_in_8_3_rest_V => fifo_in(8*NFIFOS+3).rest,
                     fifo_in_8_4_rest_V => fifo_in(8*NFIFOS+4).rest,
                     fifo_in_8_5_rest_V => fifo_in(8*NFIFOS+5).rest,
                     fifo_write_0_0 => fifo_in_write(0*NFIFOS+0),
                     fifo_write_0_1 => fifo_in_write(0*NFIFOS+1),
                     fifo_write_0_2 => fifo_in_write(0*NFIFOS+2),
                     fifo_write_0_3 => fifo_in_write(0*NFIFOS+3),
                     fifo_write_0_4 => fifo_in_write(0*NFIFOS+4),
                     fifo_write_0_5 => fifo_in_write(0*NFIFOS+5),
                     fifo_write_1_0 => fifo_in_write(1*NFIFOS+0),
                     fifo_write_1_1 => fifo_in_write(1*NFIFOS+1),
                     fifo_write_1_2 => fifo_in_write(1*NFIFOS+2),
                     fifo_write_1_3 => fifo_in_write(1*NFIFOS+3),
                     fifo_write_1_4 => fifo_in_write(1*NFIFOS+4),
                     fifo_write_1_5 => fifo_in_write(1*NFIFOS+5),
                     fifo_write_2_0 => fifo_in_write(2*NFIFOS+0),
                     fifo_write_2_1 => fifo_in_write(2*NFIFOS+1),
                     fifo_write_2_2 => fifo_in_write(2*NFIFOS+2),
                     fifo_write_2_3 => fifo_in_write(2*NFIFOS+3),
                     fifo_write_2_4 => fifo_in_write(2*NFIFOS+4),
                     fifo_write_2_5 => fifo_in_write(2*NFIFOS+5),
                     fifo_write_3_0 => fifo_in_write(3*NFIFOS+0),
                     fifo_write_3_1 => fifo_in_write(3*NFIFOS+1),
                     fifo_write_3_2 => fifo_in_write(3*NFIFOS+2),
                     fifo_write_3_3 => fifo_in_write(3*NFIFOS+3),
                     fifo_write_3_4 => fifo_in_write(3*NFIFOS+4),
                     fifo_write_3_5 => fifo_in_write(3*NFIFOS+5),
                     fifo_write_4_0 => fifo_in_write(4*NFIFOS+0),
                     fifo_write_4_1 => fifo_in_write(4*NFIFOS+1),
                     fifo_write_4_2 => fifo_in_write(4*NFIFOS+2),
                     fifo_write_4_3 => fifo_in_write(4*NFIFOS+3),
                     fifo_write_4_4 => fifo_in_write(4*NFIFOS+4),
                     fifo_write_4_5 => fifo_in_write(4*NFIFOS+5),
                     fifo_write_5_0 => fifo_in_write(5*NFIFOS+0),
                     fifo_write_5_1 => fifo_in_write(5*NFIFOS+1),
                     fifo_write_5_2 => fifo_in_write(5*NFIFOS+2),
                     fifo_write_5_3 => fifo_in_write(5*NFIFOS+3),
                     fifo_write_5_4 => fifo_in_write(5*NFIFOS+4),
                     fifo_write_5_5 => fifo_in_write(5*NFIFOS+5),
                     fifo_write_6_0 => fifo_in_write(6*NFIFOS+0),
                     fifo_write_6_1 => fifo_in_write(6*NFIFOS+1),
                     fifo_write_6_2 => fifo_in_write(6*NFIFOS+2),
                     fifo_write_6_3 => fifo_in_write(6*NFIFOS+3),
                     fifo_write_6_4 => fifo_in_write(6*NFIFOS+4),
                     fifo_write_6_5 => fifo_in_write(6*NFIFOS+5),
                     fifo_write_7_0 => fifo_in_write(7*NFIFOS+0),
                     fifo_write_7_1 => fifo_in_write(7*NFIFOS+1),
                     fifo_write_7_2 => fifo_in_write(7*NFIFOS+2),
                     fifo_write_7_3 => fifo_in_write(7*NFIFOS+3),
                     fifo_write_7_4 => fifo_in_write(7*NFIFOS+4),
                     fifo_write_7_5 => fifo_in_write(7*NFIFOS+5),
                     fifo_write_8_0 => fifo_in_write(8*NFIFOS+0),
                     fifo_write_8_1 => fifo_in_write(8*NFIFOS+1),
                     fifo_write_8_2 => fifo_in_write(8*NFIFOS+2),
                     fifo_write_8_3 => fifo_in_write(8*NFIFOS+3),
                     fifo_write_8_4 => fifo_in_write(8*NFIFOS+4),
                     fifo_write_8_5 => fifo_in_write(8*NFIFOS+5),
                     fifo_out_0_0_pt_V => fifo_out(0*NFIFOS+0).pt,
                     fifo_out_0_1_pt_V => fifo_out(0*NFIFOS+1).pt,
                     fifo_out_0_2_pt_V => fifo_out(0*NFIFOS+2).pt,
                     fifo_out_0_3_pt_V => fifo_out(0*NFIFOS+3).pt,
                     fifo_out_0_4_pt_V => fifo_out(0*NFIFOS+4).pt,
                     fifo_out_0_5_pt_V => fifo_out(0*NFIFOS+5).pt,
                     fifo_out_0_0_eta_V => fifo_out(0*NFIFOS+0).eta,
                     fifo_out_0_1_eta_V => fifo_out(0*NFIFOS+1).eta,
                     fifo_out_0_2_eta_V => fifo_out(0*NFIFOS+2).eta,
                     fifo_out_0_3_eta_V => fifo_out(0*NFIFOS+3).eta,
                     fifo_out_0_4_eta_V => fifo_out(0*NFIFOS+4).eta,
                     fifo_out_0_5_eta_V => fifo_out(0*NFIFOS+5).eta,
                     fifo_out_0_0_phi_V => fifo_out(0*NFIFOS+0).phi,
                     fifo_out_0_1_phi_V => fifo_out(0*NFIFOS+1).phi,
                     fifo_out_0_2_phi_V => fifo_out(0*NFIFOS+2).phi,
                     fifo_out_0_3_phi_V => fifo_out(0*NFIFOS+3).phi,
                     fifo_out_0_4_phi_V => fifo_out(0*NFIFOS+4).phi,
                     fifo_out_0_5_phi_V => fifo_out(0*NFIFOS+5).phi,
                     fifo_out_0_0_rest_V => fifo_out(0*NFIFOS+0).rest,
                     fifo_out_0_1_rest_V => fifo_out(0*NFIFOS+1).rest,
                     fifo_out_0_2_rest_V => fifo_out(0*NFIFOS+2).rest,
                     fifo_out_0_3_rest_V => fifo_out(0*NFIFOS+3).rest,
                     fifo_out_0_4_rest_V => fifo_out(0*NFIFOS+4).rest,
                     fifo_out_0_5_rest_V => fifo_out(0*NFIFOS+5).rest,
                     fifo_out_1_0_pt_V => fifo_out(1*NFIFOS+0).pt,
                     fifo_out_1_1_pt_V => fifo_out(1*NFIFOS+1).pt,
                     fifo_out_1_2_pt_V => fifo_out(1*NFIFOS+2).pt,
                     fifo_out_1_3_pt_V => fifo_out(1*NFIFOS+3).pt,
                     fifo_out_1_4_pt_V => fifo_out(1*NFIFOS+4).pt,
                     fifo_out_1_5_pt_V => fifo_out(1*NFIFOS+5).pt,
                     fifo_out_1_0_eta_V => fifo_out(1*NFIFOS+0).eta,
                     fifo_out_1_1_eta_V => fifo_out(1*NFIFOS+1).eta,
                     fifo_out_1_2_eta_V => fifo_out(1*NFIFOS+2).eta,
                     fifo_out_1_3_eta_V => fifo_out(1*NFIFOS+3).eta,
                     fifo_out_1_4_eta_V => fifo_out(1*NFIFOS+4).eta,
                     fifo_out_1_5_eta_V => fifo_out(1*NFIFOS+5).eta,
                     fifo_out_1_0_phi_V => fifo_out(1*NFIFOS+0).phi,
                     fifo_out_1_1_phi_V => fifo_out(1*NFIFOS+1).phi,
                     fifo_out_1_2_phi_V => fifo_out(1*NFIFOS+2).phi,
                     fifo_out_1_3_phi_V => fifo_out(1*NFIFOS+3).phi,
                     fifo_out_1_4_phi_V => fifo_out(1*NFIFOS+4).phi,
                     fifo_out_1_5_phi_V => fifo_out(1*NFIFOS+5).phi,
                     fifo_out_1_0_rest_V => fifo_out(1*NFIFOS+0).rest,
                     fifo_out_1_1_rest_V => fifo_out(1*NFIFOS+1).rest,
                     fifo_out_1_2_rest_V => fifo_out(1*NFIFOS+2).rest,
                     fifo_out_1_3_rest_V => fifo_out(1*NFIFOS+3).rest,
                     fifo_out_1_4_rest_V => fifo_out(1*NFIFOS+4).rest,
                     fifo_out_1_5_rest_V => fifo_out(1*NFIFOS+5).rest,
                     fifo_out_2_0_pt_V => fifo_out(2*NFIFOS+0).pt,
                     fifo_out_2_1_pt_V => fifo_out(2*NFIFOS+1).pt,
                     fifo_out_2_2_pt_V => fifo_out(2*NFIFOS+2).pt,
                     fifo_out_2_3_pt_V => fifo_out(2*NFIFOS+3).pt,
                     fifo_out_2_4_pt_V => fifo_out(2*NFIFOS+4).pt,
                     fifo_out_2_5_pt_V => fifo_out(2*NFIFOS+5).pt,
                     fifo_out_2_0_eta_V => fifo_out(2*NFIFOS+0).eta,
                     fifo_out_2_1_eta_V => fifo_out(2*NFIFOS+1).eta,
                     fifo_out_2_2_eta_V => fifo_out(2*NFIFOS+2).eta,
                     fifo_out_2_3_eta_V => fifo_out(2*NFIFOS+3).eta,
                     fifo_out_2_4_eta_V => fifo_out(2*NFIFOS+4).eta,
                     fifo_out_2_5_eta_V => fifo_out(2*NFIFOS+5).eta,
                     fifo_out_2_0_phi_V => fifo_out(2*NFIFOS+0).phi,
                     fifo_out_2_1_phi_V => fifo_out(2*NFIFOS+1).phi,
                     fifo_out_2_2_phi_V => fifo_out(2*NFIFOS+2).phi,
                     fifo_out_2_3_phi_V => fifo_out(2*NFIFOS+3).phi,
                     fifo_out_2_4_phi_V => fifo_out(2*NFIFOS+4).phi,
                     fifo_out_2_5_phi_V => fifo_out(2*NFIFOS+5).phi,
                     fifo_out_2_0_rest_V => fifo_out(2*NFIFOS+0).rest,
                     fifo_out_2_1_rest_V => fifo_out(2*NFIFOS+1).rest,
                     fifo_out_2_2_rest_V => fifo_out(2*NFIFOS+2).rest,
                     fifo_out_2_3_rest_V => fifo_out(2*NFIFOS+3).rest,
                     fifo_out_2_4_rest_V => fifo_out(2*NFIFOS+4).rest,
                     fifo_out_2_5_rest_V => fifo_out(2*NFIFOS+5).rest,
                     fifo_out_3_0_pt_V => fifo_out(3*NFIFOS+0).pt,
                     fifo_out_3_1_pt_V => fifo_out(3*NFIFOS+1).pt,
                     fifo_out_3_2_pt_V => fifo_out(3*NFIFOS+2).pt,
                     fifo_out_3_3_pt_V => fifo_out(3*NFIFOS+3).pt,
                     fifo_out_3_4_pt_V => fifo_out(3*NFIFOS+4).pt,
                     fifo_out_3_5_pt_V => fifo_out(3*NFIFOS+5).pt,
                     fifo_out_3_0_eta_V => fifo_out(3*NFIFOS+0).eta,
                     fifo_out_3_1_eta_V => fifo_out(3*NFIFOS+1).eta,
                     fifo_out_3_2_eta_V => fifo_out(3*NFIFOS+2).eta,
                     fifo_out_3_3_eta_V => fifo_out(3*NFIFOS+3).eta,
                     fifo_out_3_4_eta_V => fifo_out(3*NFIFOS+4).eta,
                     fifo_out_3_5_eta_V => fifo_out(3*NFIFOS+5).eta,
                     fifo_out_3_0_phi_V => fifo_out(3*NFIFOS+0).phi,
                     fifo_out_3_1_phi_V => fifo_out(3*NFIFOS+1).phi,
                     fifo_out_3_2_phi_V => fifo_out(3*NFIFOS+2).phi,
                     fifo_out_3_3_phi_V => fifo_out(3*NFIFOS+3).phi,
                     fifo_out_3_4_phi_V => fifo_out(3*NFIFOS+4).phi,
                     fifo_out_3_5_phi_V => fifo_out(3*NFIFOS+5).phi,
                     fifo_out_3_0_rest_V => fifo_out(3*NFIFOS+0).rest,
                     fifo_out_3_1_rest_V => fifo_out(3*NFIFOS+1).rest,
                     fifo_out_3_2_rest_V => fifo_out(3*NFIFOS+2).rest,
                     fifo_out_3_3_rest_V => fifo_out(3*NFIFOS+3).rest,
                     fifo_out_3_4_rest_V => fifo_out(3*NFIFOS+4).rest,
                     fifo_out_3_5_rest_V => fifo_out(3*NFIFOS+5).rest,
                     fifo_out_4_0_pt_V => fifo_out(4*NFIFOS+0).pt,
                     fifo_out_4_1_pt_V => fifo_out(4*NFIFOS+1).pt,
                     fifo_out_4_2_pt_V => fifo_out(4*NFIFOS+2).pt,
                     fifo_out_4_3_pt_V => fifo_out(4*NFIFOS+3).pt,
                     fifo_out_4_4_pt_V => fifo_out(4*NFIFOS+4).pt,
                     fifo_out_4_5_pt_V => fifo_out(4*NFIFOS+5).pt,
                     fifo_out_4_0_eta_V => fifo_out(4*NFIFOS+0).eta,
                     fifo_out_4_1_eta_V => fifo_out(4*NFIFOS+1).eta,
                     fifo_out_4_2_eta_V => fifo_out(4*NFIFOS+2).eta,
                     fifo_out_4_3_eta_V => fifo_out(4*NFIFOS+3).eta,
                     fifo_out_4_4_eta_V => fifo_out(4*NFIFOS+4).eta,
                     fifo_out_4_5_eta_V => fifo_out(4*NFIFOS+5).eta,
                     fifo_out_4_0_phi_V => fifo_out(4*NFIFOS+0).phi,
                     fifo_out_4_1_phi_V => fifo_out(4*NFIFOS+1).phi,
                     fifo_out_4_2_phi_V => fifo_out(4*NFIFOS+2).phi,
                     fifo_out_4_3_phi_V => fifo_out(4*NFIFOS+3).phi,
                     fifo_out_4_4_phi_V => fifo_out(4*NFIFOS+4).phi,
                     fifo_out_4_5_phi_V => fifo_out(4*NFIFOS+5).phi,
                     fifo_out_4_0_rest_V => fifo_out(4*NFIFOS+0).rest,
                     fifo_out_4_1_rest_V => fifo_out(4*NFIFOS+1).rest,
                     fifo_out_4_2_rest_V => fifo_out(4*NFIFOS+2).rest,
                     fifo_out_4_3_rest_V => fifo_out(4*NFIFOS+3).rest,
                     fifo_out_4_4_rest_V => fifo_out(4*NFIFOS+4).rest,
                     fifo_out_4_5_rest_V => fifo_out(4*NFIFOS+5).rest,
                     fifo_out_5_0_pt_V => fifo_out(5*NFIFOS+0).pt,
                     fifo_out_5_1_pt_V => fifo_out(5*NFIFOS+1).pt,
                     fifo_out_5_2_pt_V => fifo_out(5*NFIFOS+2).pt,
                     fifo_out_5_3_pt_V => fifo_out(5*NFIFOS+3).pt,
                     fifo_out_5_4_pt_V => fifo_out(5*NFIFOS+4).pt,
                     fifo_out_5_5_pt_V => fifo_out(5*NFIFOS+5).pt,
                     fifo_out_5_0_eta_V => fifo_out(5*NFIFOS+0).eta,
                     fifo_out_5_1_eta_V => fifo_out(5*NFIFOS+1).eta,
                     fifo_out_5_2_eta_V => fifo_out(5*NFIFOS+2).eta,
                     fifo_out_5_3_eta_V => fifo_out(5*NFIFOS+3).eta,
                     fifo_out_5_4_eta_V => fifo_out(5*NFIFOS+4).eta,
                     fifo_out_5_5_eta_V => fifo_out(5*NFIFOS+5).eta,
                     fifo_out_5_0_phi_V => fifo_out(5*NFIFOS+0).phi,
                     fifo_out_5_1_phi_V => fifo_out(5*NFIFOS+1).phi,
                     fifo_out_5_2_phi_V => fifo_out(5*NFIFOS+2).phi,
                     fifo_out_5_3_phi_V => fifo_out(5*NFIFOS+3).phi,
                     fifo_out_5_4_phi_V => fifo_out(5*NFIFOS+4).phi,
                     fifo_out_5_5_phi_V => fifo_out(5*NFIFOS+5).phi,
                     fifo_out_5_0_rest_V => fifo_out(5*NFIFOS+0).rest,
                     fifo_out_5_1_rest_V => fifo_out(5*NFIFOS+1).rest,
                     fifo_out_5_2_rest_V => fifo_out(5*NFIFOS+2).rest,
                     fifo_out_5_3_rest_V => fifo_out(5*NFIFOS+3).rest,
                     fifo_out_5_4_rest_V => fifo_out(5*NFIFOS+4).rest,
                     fifo_out_5_5_rest_V => fifo_out(5*NFIFOS+5).rest,
                     fifo_out_6_0_pt_V => fifo_out(6*NFIFOS+0).pt,
                     fifo_out_6_1_pt_V => fifo_out(6*NFIFOS+1).pt,
                     fifo_out_6_2_pt_V => fifo_out(6*NFIFOS+2).pt,
                     fifo_out_6_3_pt_V => fifo_out(6*NFIFOS+3).pt,
                     fifo_out_6_4_pt_V => fifo_out(6*NFIFOS+4).pt,
                     fifo_out_6_5_pt_V => fifo_out(6*NFIFOS+5).pt,
                     fifo_out_6_0_eta_V => fifo_out(6*NFIFOS+0).eta,
                     fifo_out_6_1_eta_V => fifo_out(6*NFIFOS+1).eta,
                     fifo_out_6_2_eta_V => fifo_out(6*NFIFOS+2).eta,
                     fifo_out_6_3_eta_V => fifo_out(6*NFIFOS+3).eta,
                     fifo_out_6_4_eta_V => fifo_out(6*NFIFOS+4).eta,
                     fifo_out_6_5_eta_V => fifo_out(6*NFIFOS+5).eta,
                     fifo_out_6_0_phi_V => fifo_out(6*NFIFOS+0).phi,
                     fifo_out_6_1_phi_V => fifo_out(6*NFIFOS+1).phi,
                     fifo_out_6_2_phi_V => fifo_out(6*NFIFOS+2).phi,
                     fifo_out_6_3_phi_V => fifo_out(6*NFIFOS+3).phi,
                     fifo_out_6_4_phi_V => fifo_out(6*NFIFOS+4).phi,
                     fifo_out_6_5_phi_V => fifo_out(6*NFIFOS+5).phi,
                     fifo_out_6_0_rest_V => fifo_out(6*NFIFOS+0).rest,
                     fifo_out_6_1_rest_V => fifo_out(6*NFIFOS+1).rest,
                     fifo_out_6_2_rest_V => fifo_out(6*NFIFOS+2).rest,
                     fifo_out_6_3_rest_V => fifo_out(6*NFIFOS+3).rest,
                     fifo_out_6_4_rest_V => fifo_out(6*NFIFOS+4).rest,
                     fifo_out_6_5_rest_V => fifo_out(6*NFIFOS+5).rest,
                     fifo_out_7_0_pt_V => fifo_out(7*NFIFOS+0).pt,
                     fifo_out_7_1_pt_V => fifo_out(7*NFIFOS+1).pt,
                     fifo_out_7_2_pt_V => fifo_out(7*NFIFOS+2).pt,
                     fifo_out_7_3_pt_V => fifo_out(7*NFIFOS+3).pt,
                     fifo_out_7_4_pt_V => fifo_out(7*NFIFOS+4).pt,
                     fifo_out_7_5_pt_V => fifo_out(7*NFIFOS+5).pt,
                     fifo_out_7_0_eta_V => fifo_out(7*NFIFOS+0).eta,
                     fifo_out_7_1_eta_V => fifo_out(7*NFIFOS+1).eta,
                     fifo_out_7_2_eta_V => fifo_out(7*NFIFOS+2).eta,
                     fifo_out_7_3_eta_V => fifo_out(7*NFIFOS+3).eta,
                     fifo_out_7_4_eta_V => fifo_out(7*NFIFOS+4).eta,
                     fifo_out_7_5_eta_V => fifo_out(7*NFIFOS+5).eta,
                     fifo_out_7_0_phi_V => fifo_out(7*NFIFOS+0).phi,
                     fifo_out_7_1_phi_V => fifo_out(7*NFIFOS+1).phi,
                     fifo_out_7_2_phi_V => fifo_out(7*NFIFOS+2).phi,
                     fifo_out_7_3_phi_V => fifo_out(7*NFIFOS+3).phi,
                     fifo_out_7_4_phi_V => fifo_out(7*NFIFOS+4).phi,
                     fifo_out_7_5_phi_V => fifo_out(7*NFIFOS+5).phi,
                     fifo_out_7_0_rest_V => fifo_out(7*NFIFOS+0).rest,
                     fifo_out_7_1_rest_V => fifo_out(7*NFIFOS+1).rest,
                     fifo_out_7_2_rest_V => fifo_out(7*NFIFOS+2).rest,
                     fifo_out_7_3_rest_V => fifo_out(7*NFIFOS+3).rest,
                     fifo_out_7_4_rest_V => fifo_out(7*NFIFOS+4).rest,
                     fifo_out_7_5_rest_V => fifo_out(7*NFIFOS+5).rest,
                     fifo_out_8_0_pt_V => fifo_out(8*NFIFOS+0).pt,
                     fifo_out_8_1_pt_V => fifo_out(8*NFIFOS+1).pt,
                     fifo_out_8_2_pt_V => fifo_out(8*NFIFOS+2).pt,
                     fifo_out_8_3_pt_V => fifo_out(8*NFIFOS+3).pt,
                     fifo_out_8_4_pt_V => fifo_out(8*NFIFOS+4).pt,
                     fifo_out_8_5_pt_V => fifo_out(8*NFIFOS+5).pt,
                     fifo_out_8_0_eta_V => fifo_out(8*NFIFOS+0).eta,
                     fifo_out_8_1_eta_V => fifo_out(8*NFIFOS+1).eta,
                     fifo_out_8_2_eta_V => fifo_out(8*NFIFOS+2).eta,
                     fifo_out_8_3_eta_V => fifo_out(8*NFIFOS+3).eta,
                     fifo_out_8_4_eta_V => fifo_out(8*NFIFOS+4).eta,
                     fifo_out_8_5_eta_V => fifo_out(8*NFIFOS+5).eta,
                     fifo_out_8_0_phi_V => fifo_out(8*NFIFOS+0).phi,
                     fifo_out_8_1_phi_V => fifo_out(8*NFIFOS+1).phi,
                     fifo_out_8_2_phi_V => fifo_out(8*NFIFOS+2).phi,
                     fifo_out_8_3_phi_V => fifo_out(8*NFIFOS+3).phi,
                     fifo_out_8_4_phi_V => fifo_out(8*NFIFOS+4).phi,
                     fifo_out_8_5_phi_V => fifo_out(8*NFIFOS+5).phi,
                     fifo_out_8_0_rest_V => fifo_out(8*NFIFOS+0).rest,
                     fifo_out_8_1_rest_V => fifo_out(8*NFIFOS+1).rest,
                     fifo_out_8_2_rest_V => fifo_out(8*NFIFOS+2).rest,
                     fifo_out_8_3_rest_V => fifo_out(8*NFIFOS+3).rest,
                     fifo_out_8_4_rest_V => fifo_out(8*NFIFOS+4).rest,
                     fifo_out_8_5_rest_V => fifo_out(8*NFIFOS+5).rest,
                     fifo_out_valid_0_0 => fifo_out_valid(0*NFIFOS+0),
                     fifo_out_valid_0_1 => fifo_out_valid(0*NFIFOS+1),
                     fifo_out_valid_0_2 => fifo_out_valid(0*NFIFOS+2),
                     fifo_out_valid_0_3 => fifo_out_valid(0*NFIFOS+3),
                     fifo_out_valid_0_4 => fifo_out_valid(0*NFIFOS+4),
                     fifo_out_valid_0_5 => fifo_out_valid(0*NFIFOS+5),
                     fifo_out_valid_1_0 => fifo_out_valid(1*NFIFOS+0),
                     fifo_out_valid_1_1 => fifo_out_valid(1*NFIFOS+1),
                     fifo_out_valid_1_2 => fifo_out_valid(1*NFIFOS+2),
                     fifo_out_valid_1_3 => fifo_out_valid(1*NFIFOS+3),
                     fifo_out_valid_1_4 => fifo_out_valid(1*NFIFOS+4),
                     fifo_out_valid_1_5 => fifo_out_valid(1*NFIFOS+5),
                     fifo_out_valid_2_0 => fifo_out_valid(2*NFIFOS+0),
                     fifo_out_valid_2_1 => fifo_out_valid(2*NFIFOS+1),
                     fifo_out_valid_2_2 => fifo_out_valid(2*NFIFOS+2),
                     fifo_out_valid_2_3 => fifo_out_valid(2*NFIFOS+3),
                     fifo_out_valid_2_4 => fifo_out_valid(2*NFIFOS+4),
                     fifo_out_valid_2_5 => fifo_out_valid(2*NFIFOS+5),
                     fifo_out_valid_3_0 => fifo_out_valid(3*NFIFOS+0),
                     fifo_out_valid_3_1 => fifo_out_valid(3*NFIFOS+1),
                     fifo_out_valid_3_2 => fifo_out_valid(3*NFIFOS+2),
                     fifo_out_valid_3_3 => fifo_out_valid(3*NFIFOS+3),
                     fifo_out_valid_3_4 => fifo_out_valid(3*NFIFOS+4),
                     fifo_out_valid_3_5 => fifo_out_valid(3*NFIFOS+5),
                     fifo_out_valid_4_0 => fifo_out_valid(4*NFIFOS+0),
                     fifo_out_valid_4_1 => fifo_out_valid(4*NFIFOS+1),
                     fifo_out_valid_4_2 => fifo_out_valid(4*NFIFOS+2),
                     fifo_out_valid_4_3 => fifo_out_valid(4*NFIFOS+3),
                     fifo_out_valid_4_4 => fifo_out_valid(4*NFIFOS+4),
                     fifo_out_valid_4_5 => fifo_out_valid(4*NFIFOS+5),
                     fifo_out_valid_5_0 => fifo_out_valid(5*NFIFOS+0),
                     fifo_out_valid_5_1 => fifo_out_valid(5*NFIFOS+1),
                     fifo_out_valid_5_2 => fifo_out_valid(5*NFIFOS+2),
                     fifo_out_valid_5_3 => fifo_out_valid(5*NFIFOS+3),
                     fifo_out_valid_5_4 => fifo_out_valid(5*NFIFOS+4),
                     fifo_out_valid_5_5 => fifo_out_valid(5*NFIFOS+5),
                     fifo_out_valid_6_0 => fifo_out_valid(6*NFIFOS+0),
                     fifo_out_valid_6_1 => fifo_out_valid(6*NFIFOS+1),
                     fifo_out_valid_6_2 => fifo_out_valid(6*NFIFOS+2),
                     fifo_out_valid_6_3 => fifo_out_valid(6*NFIFOS+3),
                     fifo_out_valid_6_4 => fifo_out_valid(6*NFIFOS+4),
                     fifo_out_valid_6_5 => fifo_out_valid(6*NFIFOS+5),
                     fifo_out_valid_7_0 => fifo_out_valid(7*NFIFOS+0),
                     fifo_out_valid_7_1 => fifo_out_valid(7*NFIFOS+1),
                     fifo_out_valid_7_2 => fifo_out_valid(7*NFIFOS+2),
                     fifo_out_valid_7_3 => fifo_out_valid(7*NFIFOS+3),
                     fifo_out_valid_7_4 => fifo_out_valid(7*NFIFOS+4),
                     fifo_out_valid_7_5 => fifo_out_valid(7*NFIFOS+5),
                     fifo_out_valid_8_0 => fifo_out_valid(8*NFIFOS+0),
                     fifo_out_valid_8_1 => fifo_out_valid(8*NFIFOS+1),
                     fifo_out_valid_8_2 => fifo_out_valid(8*NFIFOS+2),
                     fifo_out_valid_8_3 => fifo_out_valid(8*NFIFOS+3),
                     fifo_out_valid_8_4 => fifo_out_valid(8*NFIFOS+4),
                     fifo_out_valid_8_5 => fifo_out_valid(8*NFIFOS+5),
                     fifo_out_roll_0_0 => fifo_out_roll(0*NFIFOS+0),
                     fifo_out_roll_0_1 => fifo_out_roll(0*NFIFOS+1),
                     fifo_out_roll_0_2 => fifo_out_roll(0*NFIFOS+2),
                     fifo_out_roll_0_3 => fifo_out_roll(0*NFIFOS+3),
                     fifo_out_roll_0_4 => fifo_out_roll(0*NFIFOS+4),
                     fifo_out_roll_0_5 => fifo_out_roll(0*NFIFOS+5),
                     fifo_out_roll_1_0 => fifo_out_roll(1*NFIFOS+0),
                     fifo_out_roll_1_1 => fifo_out_roll(1*NFIFOS+1),
                     fifo_out_roll_1_2 => fifo_out_roll(1*NFIFOS+2),
                     fifo_out_roll_1_3 => fifo_out_roll(1*NFIFOS+3),
                     fifo_out_roll_1_4 => fifo_out_roll(1*NFIFOS+4),
                     fifo_out_roll_1_5 => fifo_out_roll(1*NFIFOS+5),
                     fifo_out_roll_2_0 => fifo_out_roll(2*NFIFOS+0),
                     fifo_out_roll_2_1 => fifo_out_roll(2*NFIFOS+1),
                     fifo_out_roll_2_2 => fifo_out_roll(2*NFIFOS+2),
                     fifo_out_roll_2_3 => fifo_out_roll(2*NFIFOS+3),
                     fifo_out_roll_2_4 => fifo_out_roll(2*NFIFOS+4),
                     fifo_out_roll_2_5 => fifo_out_roll(2*NFIFOS+5),
                     fifo_out_roll_3_0 => fifo_out_roll(3*NFIFOS+0),
                     fifo_out_roll_3_1 => fifo_out_roll(3*NFIFOS+1),
                     fifo_out_roll_3_2 => fifo_out_roll(3*NFIFOS+2),
                     fifo_out_roll_3_3 => fifo_out_roll(3*NFIFOS+3),
                     fifo_out_roll_3_4 => fifo_out_roll(3*NFIFOS+4),
                     fifo_out_roll_3_5 => fifo_out_roll(3*NFIFOS+5),
                     fifo_out_roll_4_0 => fifo_out_roll(4*NFIFOS+0),
                     fifo_out_roll_4_1 => fifo_out_roll(4*NFIFOS+1),
                     fifo_out_roll_4_2 => fifo_out_roll(4*NFIFOS+2),
                     fifo_out_roll_4_3 => fifo_out_roll(4*NFIFOS+3),
                     fifo_out_roll_4_4 => fifo_out_roll(4*NFIFOS+4),
                     fifo_out_roll_4_5 => fifo_out_roll(4*NFIFOS+5),
                     fifo_out_roll_5_0 => fifo_out_roll(5*NFIFOS+0),
                     fifo_out_roll_5_1 => fifo_out_roll(5*NFIFOS+1),
                     fifo_out_roll_5_2 => fifo_out_roll(5*NFIFOS+2),
                     fifo_out_roll_5_3 => fifo_out_roll(5*NFIFOS+3),
                     fifo_out_roll_5_4 => fifo_out_roll(5*NFIFOS+4),
                     fifo_out_roll_5_5 => fifo_out_roll(5*NFIFOS+5),
                     fifo_out_roll_6_0 => fifo_out_roll(6*NFIFOS+0),
                     fifo_out_roll_6_1 => fifo_out_roll(6*NFIFOS+1),
                     fifo_out_roll_6_2 => fifo_out_roll(6*NFIFOS+2),
                     fifo_out_roll_6_3 => fifo_out_roll(6*NFIFOS+3),
                     fifo_out_roll_6_4 => fifo_out_roll(6*NFIFOS+4),
                     fifo_out_roll_6_5 => fifo_out_roll(6*NFIFOS+5),
                     fifo_out_roll_7_0 => fifo_out_roll(7*NFIFOS+0),
                     fifo_out_roll_7_1 => fifo_out_roll(7*NFIFOS+1),
                     fifo_out_roll_7_2 => fifo_out_roll(7*NFIFOS+2),
                     fifo_out_roll_7_3 => fifo_out_roll(7*NFIFOS+3),
                     fifo_out_roll_7_4 => fifo_out_roll(7*NFIFOS+4),
                     fifo_out_roll_7_5 => fifo_out_roll(7*NFIFOS+5),
                     fifo_out_roll_8_0 => fifo_out_roll(8*NFIFOS+0),
                     fifo_out_roll_8_1 => fifo_out_roll(8*NFIFOS+1),
                     fifo_out_roll_8_2 => fifo_out_roll(8*NFIFOS+2),
                     fifo_out_roll_8_3 => fifo_out_roll(8*NFIFOS+3),
                     fifo_out_roll_8_4 => fifo_out_roll(8*NFIFOS+4),
                     fifo_out_roll_8_5 => fifo_out_roll(8*NFIFOS+5),
                     fifo_full_0_0 => fifo_out_full(0*NFIFOS+0),
                     fifo_full_0_1 => fifo_out_full(0*NFIFOS+1),
                     fifo_full_0_2 => fifo_out_full(0*NFIFOS+2),
                     fifo_full_0_3 => fifo_out_full(0*NFIFOS+3),
                     fifo_full_0_4 => fifo_out_full(0*NFIFOS+4),
                     fifo_full_0_5 => fifo_out_full(0*NFIFOS+5),
                     fifo_full_1_0 => fifo_out_full(1*NFIFOS+0),
                     fifo_full_1_1 => fifo_out_full(1*NFIFOS+1),
                     fifo_full_1_2 => fifo_out_full(1*NFIFOS+2),
                     fifo_full_1_3 => fifo_out_full(1*NFIFOS+3),
                     fifo_full_1_4 => fifo_out_full(1*NFIFOS+4),
                     fifo_full_1_5 => fifo_out_full(1*NFIFOS+5),
                     fifo_full_2_0 => fifo_out_full(2*NFIFOS+0),
                     fifo_full_2_1 => fifo_out_full(2*NFIFOS+1),
                     fifo_full_2_2 => fifo_out_full(2*NFIFOS+2),
                     fifo_full_2_3 => fifo_out_full(2*NFIFOS+3),
                     fifo_full_2_4 => fifo_out_full(2*NFIFOS+4),
                     fifo_full_2_5 => fifo_out_full(2*NFIFOS+5),
                     fifo_full_3_0 => fifo_out_full(3*NFIFOS+0),
                     fifo_full_3_1 => fifo_out_full(3*NFIFOS+1),
                     fifo_full_3_2 => fifo_out_full(3*NFIFOS+2),
                     fifo_full_3_3 => fifo_out_full(3*NFIFOS+3),
                     fifo_full_3_4 => fifo_out_full(3*NFIFOS+4),
                     fifo_full_3_5 => fifo_out_full(3*NFIFOS+5),
                     fifo_full_4_0 => fifo_out_full(4*NFIFOS+0),
                     fifo_full_4_1 => fifo_out_full(4*NFIFOS+1),
                     fifo_full_4_2 => fifo_out_full(4*NFIFOS+2),
                     fifo_full_4_3 => fifo_out_full(4*NFIFOS+3),
                     fifo_full_4_4 => fifo_out_full(4*NFIFOS+4),
                     fifo_full_4_5 => fifo_out_full(4*NFIFOS+5),
                     fifo_full_5_0 => fifo_out_full(5*NFIFOS+0),
                     fifo_full_5_1 => fifo_out_full(5*NFIFOS+1),
                     fifo_full_5_2 => fifo_out_full(5*NFIFOS+2),
                     fifo_full_5_3 => fifo_out_full(5*NFIFOS+3),
                     fifo_full_5_4 => fifo_out_full(5*NFIFOS+4),
                     fifo_full_5_5 => fifo_out_full(5*NFIFOS+5),
                     fifo_full_6_0 => fifo_out_full(6*NFIFOS+0),
                     fifo_full_6_1 => fifo_out_full(6*NFIFOS+1),
                     fifo_full_6_2 => fifo_out_full(6*NFIFOS+2),
                     fifo_full_6_3 => fifo_out_full(6*NFIFOS+3),
                     fifo_full_6_4 => fifo_out_full(6*NFIFOS+4),
                     fifo_full_6_5 => fifo_out_full(6*NFIFOS+5),
                     fifo_full_7_0 => fifo_out_full(7*NFIFOS+0),
                     fifo_full_7_1 => fifo_out_full(7*NFIFOS+1),
                     fifo_full_7_2 => fifo_out_full(7*NFIFOS+2),
                     fifo_full_7_3 => fifo_out_full(7*NFIFOS+3),
                     fifo_full_7_4 => fifo_out_full(7*NFIFOS+4),
                     fifo_full_7_5 => fifo_out_full(7*NFIFOS+5),
                     fifo_full_8_0 => fifo_out_full(8*NFIFOS+0),
                     fifo_full_8_1 => fifo_out_full(8*NFIFOS+1),
                     fifo_full_8_2 => fifo_out_full(8*NFIFOS+2),
                     fifo_full_8_3 => fifo_out_full(8*NFIFOS+3),
                     fifo_full_8_4 => fifo_out_full(8*NFIFOS+4),
                     fifo_full_8_5 => fifo_out_full(8*NFIFOS+5)
                 );


    merge2_slice : entity work.router_merge2_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     fifo_out_0_0_pt_V => fifo_out(0*NFIFOS+0).pt,
                     fifo_out_0_1_pt_V => fifo_out(0*NFIFOS+1).pt,
                     fifo_out_0_2_pt_V => fifo_out(0*NFIFOS+2).pt,
                     fifo_out_0_3_pt_V => fifo_out(0*NFIFOS+3).pt,
                     fifo_out_0_4_pt_V => fifo_out(0*NFIFOS+4).pt,
                     fifo_out_0_5_pt_V => fifo_out(0*NFIFOS+5).pt,
                     fifo_out_0_0_eta_V => fifo_out(0*NFIFOS+0).eta,
                     fifo_out_0_1_eta_V => fifo_out(0*NFIFOS+1).eta,
                     fifo_out_0_2_eta_V => fifo_out(0*NFIFOS+2).eta,
                     fifo_out_0_3_eta_V => fifo_out(0*NFIFOS+3).eta,
                     fifo_out_0_4_eta_V => fifo_out(0*NFIFOS+4).eta,
                     fifo_out_0_5_eta_V => fifo_out(0*NFIFOS+5).eta,
                     fifo_out_0_0_phi_V => fifo_out(0*NFIFOS+0).phi,
                     fifo_out_0_1_phi_V => fifo_out(0*NFIFOS+1).phi,
                     fifo_out_0_2_phi_V => fifo_out(0*NFIFOS+2).phi,
                     fifo_out_0_3_phi_V => fifo_out(0*NFIFOS+3).phi,
                     fifo_out_0_4_phi_V => fifo_out(0*NFIFOS+4).phi,
                     fifo_out_0_5_phi_V => fifo_out(0*NFIFOS+5).phi,
                     fifo_out_0_0_rest_V => fifo_out(0*NFIFOS+0).rest,
                     fifo_out_0_1_rest_V => fifo_out(0*NFIFOS+1).rest,
                     fifo_out_0_2_rest_V => fifo_out(0*NFIFOS+2).rest,
                     fifo_out_0_3_rest_V => fifo_out(0*NFIFOS+3).rest,
                     fifo_out_0_4_rest_V => fifo_out(0*NFIFOS+4).rest,
                     fifo_out_0_5_rest_V => fifo_out(0*NFIFOS+5).rest,
                     fifo_out_1_0_pt_V => fifo_out(1*NFIFOS+0).pt,
                     fifo_out_1_1_pt_V => fifo_out(1*NFIFOS+1).pt,
                     fifo_out_1_2_pt_V => fifo_out(1*NFIFOS+2).pt,
                     fifo_out_1_3_pt_V => fifo_out(1*NFIFOS+3).pt,
                     fifo_out_1_4_pt_V => fifo_out(1*NFIFOS+4).pt,
                     fifo_out_1_5_pt_V => fifo_out(1*NFIFOS+5).pt,
                     fifo_out_1_0_eta_V => fifo_out(1*NFIFOS+0).eta,
                     fifo_out_1_1_eta_V => fifo_out(1*NFIFOS+1).eta,
                     fifo_out_1_2_eta_V => fifo_out(1*NFIFOS+2).eta,
                     fifo_out_1_3_eta_V => fifo_out(1*NFIFOS+3).eta,
                     fifo_out_1_4_eta_V => fifo_out(1*NFIFOS+4).eta,
                     fifo_out_1_5_eta_V => fifo_out(1*NFIFOS+5).eta,
                     fifo_out_1_0_phi_V => fifo_out(1*NFIFOS+0).phi,
                     fifo_out_1_1_phi_V => fifo_out(1*NFIFOS+1).phi,
                     fifo_out_1_2_phi_V => fifo_out(1*NFIFOS+2).phi,
                     fifo_out_1_3_phi_V => fifo_out(1*NFIFOS+3).phi,
                     fifo_out_1_4_phi_V => fifo_out(1*NFIFOS+4).phi,
                     fifo_out_1_5_phi_V => fifo_out(1*NFIFOS+5).phi,
                     fifo_out_1_0_rest_V => fifo_out(1*NFIFOS+0).rest,
                     fifo_out_1_1_rest_V => fifo_out(1*NFIFOS+1).rest,
                     fifo_out_1_2_rest_V => fifo_out(1*NFIFOS+2).rest,
                     fifo_out_1_3_rest_V => fifo_out(1*NFIFOS+3).rest,
                     fifo_out_1_4_rest_V => fifo_out(1*NFIFOS+4).rest,
                     fifo_out_1_5_rest_V => fifo_out(1*NFIFOS+5).rest,
                     fifo_out_2_0_pt_V => fifo_out(2*NFIFOS+0).pt,
                     fifo_out_2_1_pt_V => fifo_out(2*NFIFOS+1).pt,
                     fifo_out_2_2_pt_V => fifo_out(2*NFIFOS+2).pt,
                     fifo_out_2_3_pt_V => fifo_out(2*NFIFOS+3).pt,
                     fifo_out_2_4_pt_V => fifo_out(2*NFIFOS+4).pt,
                     fifo_out_2_5_pt_V => fifo_out(2*NFIFOS+5).pt,
                     fifo_out_2_0_eta_V => fifo_out(2*NFIFOS+0).eta,
                     fifo_out_2_1_eta_V => fifo_out(2*NFIFOS+1).eta,
                     fifo_out_2_2_eta_V => fifo_out(2*NFIFOS+2).eta,
                     fifo_out_2_3_eta_V => fifo_out(2*NFIFOS+3).eta,
                     fifo_out_2_4_eta_V => fifo_out(2*NFIFOS+4).eta,
                     fifo_out_2_5_eta_V => fifo_out(2*NFIFOS+5).eta,
                     fifo_out_2_0_phi_V => fifo_out(2*NFIFOS+0).phi,
                     fifo_out_2_1_phi_V => fifo_out(2*NFIFOS+1).phi,
                     fifo_out_2_2_phi_V => fifo_out(2*NFIFOS+2).phi,
                     fifo_out_2_3_phi_V => fifo_out(2*NFIFOS+3).phi,
                     fifo_out_2_4_phi_V => fifo_out(2*NFIFOS+4).phi,
                     fifo_out_2_5_phi_V => fifo_out(2*NFIFOS+5).phi,
                     fifo_out_2_0_rest_V => fifo_out(2*NFIFOS+0).rest,
                     fifo_out_2_1_rest_V => fifo_out(2*NFIFOS+1).rest,
                     fifo_out_2_2_rest_V => fifo_out(2*NFIFOS+2).rest,
                     fifo_out_2_3_rest_V => fifo_out(2*NFIFOS+3).rest,
                     fifo_out_2_4_rest_V => fifo_out(2*NFIFOS+4).rest,
                     fifo_out_2_5_rest_V => fifo_out(2*NFIFOS+5).rest,
                     fifo_out_3_0_pt_V => fifo_out(3*NFIFOS+0).pt,
                     fifo_out_3_1_pt_V => fifo_out(3*NFIFOS+1).pt,
                     fifo_out_3_2_pt_V => fifo_out(3*NFIFOS+2).pt,
                     fifo_out_3_3_pt_V => fifo_out(3*NFIFOS+3).pt,
                     fifo_out_3_4_pt_V => fifo_out(3*NFIFOS+4).pt,
                     fifo_out_3_5_pt_V => fifo_out(3*NFIFOS+5).pt,
                     fifo_out_3_0_eta_V => fifo_out(3*NFIFOS+0).eta,
                     fifo_out_3_1_eta_V => fifo_out(3*NFIFOS+1).eta,
                     fifo_out_3_2_eta_V => fifo_out(3*NFIFOS+2).eta,
                     fifo_out_3_3_eta_V => fifo_out(3*NFIFOS+3).eta,
                     fifo_out_3_4_eta_V => fifo_out(3*NFIFOS+4).eta,
                     fifo_out_3_5_eta_V => fifo_out(3*NFIFOS+5).eta,
                     fifo_out_3_0_phi_V => fifo_out(3*NFIFOS+0).phi,
                     fifo_out_3_1_phi_V => fifo_out(3*NFIFOS+1).phi,
                     fifo_out_3_2_phi_V => fifo_out(3*NFIFOS+2).phi,
                     fifo_out_3_3_phi_V => fifo_out(3*NFIFOS+3).phi,
                     fifo_out_3_4_phi_V => fifo_out(3*NFIFOS+4).phi,
                     fifo_out_3_5_phi_V => fifo_out(3*NFIFOS+5).phi,
                     fifo_out_3_0_rest_V => fifo_out(3*NFIFOS+0).rest,
                     fifo_out_3_1_rest_V => fifo_out(3*NFIFOS+1).rest,
                     fifo_out_3_2_rest_V => fifo_out(3*NFIFOS+2).rest,
                     fifo_out_3_3_rest_V => fifo_out(3*NFIFOS+3).rest,
                     fifo_out_3_4_rest_V => fifo_out(3*NFIFOS+4).rest,
                     fifo_out_3_5_rest_V => fifo_out(3*NFIFOS+5).rest,
                     fifo_out_4_0_pt_V => fifo_out(4*NFIFOS+0).pt,
                     fifo_out_4_1_pt_V => fifo_out(4*NFIFOS+1).pt,
                     fifo_out_4_2_pt_V => fifo_out(4*NFIFOS+2).pt,
                     fifo_out_4_3_pt_V => fifo_out(4*NFIFOS+3).pt,
                     fifo_out_4_4_pt_V => fifo_out(4*NFIFOS+4).pt,
                     fifo_out_4_5_pt_V => fifo_out(4*NFIFOS+5).pt,
                     fifo_out_4_0_eta_V => fifo_out(4*NFIFOS+0).eta,
                     fifo_out_4_1_eta_V => fifo_out(4*NFIFOS+1).eta,
                     fifo_out_4_2_eta_V => fifo_out(4*NFIFOS+2).eta,
                     fifo_out_4_3_eta_V => fifo_out(4*NFIFOS+3).eta,
                     fifo_out_4_4_eta_V => fifo_out(4*NFIFOS+4).eta,
                     fifo_out_4_5_eta_V => fifo_out(4*NFIFOS+5).eta,
                     fifo_out_4_0_phi_V => fifo_out(4*NFIFOS+0).phi,
                     fifo_out_4_1_phi_V => fifo_out(4*NFIFOS+1).phi,
                     fifo_out_4_2_phi_V => fifo_out(4*NFIFOS+2).phi,
                     fifo_out_4_3_phi_V => fifo_out(4*NFIFOS+3).phi,
                     fifo_out_4_4_phi_V => fifo_out(4*NFIFOS+4).phi,
                     fifo_out_4_5_phi_V => fifo_out(4*NFIFOS+5).phi,
                     fifo_out_4_0_rest_V => fifo_out(4*NFIFOS+0).rest,
                     fifo_out_4_1_rest_V => fifo_out(4*NFIFOS+1).rest,
                     fifo_out_4_2_rest_V => fifo_out(4*NFIFOS+2).rest,
                     fifo_out_4_3_rest_V => fifo_out(4*NFIFOS+3).rest,
                     fifo_out_4_4_rest_V => fifo_out(4*NFIFOS+4).rest,
                     fifo_out_4_5_rest_V => fifo_out(4*NFIFOS+5).rest,
                     fifo_out_5_0_pt_V => fifo_out(5*NFIFOS+0).pt,
                     fifo_out_5_1_pt_V => fifo_out(5*NFIFOS+1).pt,
                     fifo_out_5_2_pt_V => fifo_out(5*NFIFOS+2).pt,
                     fifo_out_5_3_pt_V => fifo_out(5*NFIFOS+3).pt,
                     fifo_out_5_4_pt_V => fifo_out(5*NFIFOS+4).pt,
                     fifo_out_5_5_pt_V => fifo_out(5*NFIFOS+5).pt,
                     fifo_out_5_0_eta_V => fifo_out(5*NFIFOS+0).eta,
                     fifo_out_5_1_eta_V => fifo_out(5*NFIFOS+1).eta,
                     fifo_out_5_2_eta_V => fifo_out(5*NFIFOS+2).eta,
                     fifo_out_5_3_eta_V => fifo_out(5*NFIFOS+3).eta,
                     fifo_out_5_4_eta_V => fifo_out(5*NFIFOS+4).eta,
                     fifo_out_5_5_eta_V => fifo_out(5*NFIFOS+5).eta,
                     fifo_out_5_0_phi_V => fifo_out(5*NFIFOS+0).phi,
                     fifo_out_5_1_phi_V => fifo_out(5*NFIFOS+1).phi,
                     fifo_out_5_2_phi_V => fifo_out(5*NFIFOS+2).phi,
                     fifo_out_5_3_phi_V => fifo_out(5*NFIFOS+3).phi,
                     fifo_out_5_4_phi_V => fifo_out(5*NFIFOS+4).phi,
                     fifo_out_5_5_phi_V => fifo_out(5*NFIFOS+5).phi,
                     fifo_out_5_0_rest_V => fifo_out(5*NFIFOS+0).rest,
                     fifo_out_5_1_rest_V => fifo_out(5*NFIFOS+1).rest,
                     fifo_out_5_2_rest_V => fifo_out(5*NFIFOS+2).rest,
                     fifo_out_5_3_rest_V => fifo_out(5*NFIFOS+3).rest,
                     fifo_out_5_4_rest_V => fifo_out(5*NFIFOS+4).rest,
                     fifo_out_5_5_rest_V => fifo_out(5*NFIFOS+5).rest,
                     fifo_out_6_0_pt_V => fifo_out(6*NFIFOS+0).pt,
                     fifo_out_6_1_pt_V => fifo_out(6*NFIFOS+1).pt,
                     fifo_out_6_2_pt_V => fifo_out(6*NFIFOS+2).pt,
                     fifo_out_6_3_pt_V => fifo_out(6*NFIFOS+3).pt,
                     fifo_out_6_4_pt_V => fifo_out(6*NFIFOS+4).pt,
                     fifo_out_6_5_pt_V => fifo_out(6*NFIFOS+5).pt,
                     fifo_out_6_0_eta_V => fifo_out(6*NFIFOS+0).eta,
                     fifo_out_6_1_eta_V => fifo_out(6*NFIFOS+1).eta,
                     fifo_out_6_2_eta_V => fifo_out(6*NFIFOS+2).eta,
                     fifo_out_6_3_eta_V => fifo_out(6*NFIFOS+3).eta,
                     fifo_out_6_4_eta_V => fifo_out(6*NFIFOS+4).eta,
                     fifo_out_6_5_eta_V => fifo_out(6*NFIFOS+5).eta,
                     fifo_out_6_0_phi_V => fifo_out(6*NFIFOS+0).phi,
                     fifo_out_6_1_phi_V => fifo_out(6*NFIFOS+1).phi,
                     fifo_out_6_2_phi_V => fifo_out(6*NFIFOS+2).phi,
                     fifo_out_6_3_phi_V => fifo_out(6*NFIFOS+3).phi,
                     fifo_out_6_4_phi_V => fifo_out(6*NFIFOS+4).phi,
                     fifo_out_6_5_phi_V => fifo_out(6*NFIFOS+5).phi,
                     fifo_out_6_0_rest_V => fifo_out(6*NFIFOS+0).rest,
                     fifo_out_6_1_rest_V => fifo_out(6*NFIFOS+1).rest,
                     fifo_out_6_2_rest_V => fifo_out(6*NFIFOS+2).rest,
                     fifo_out_6_3_rest_V => fifo_out(6*NFIFOS+3).rest,
                     fifo_out_6_4_rest_V => fifo_out(6*NFIFOS+4).rest,
                     fifo_out_6_5_rest_V => fifo_out(6*NFIFOS+5).rest,
                     fifo_out_7_0_pt_V => fifo_out(7*NFIFOS+0).pt,
                     fifo_out_7_1_pt_V => fifo_out(7*NFIFOS+1).pt,
                     fifo_out_7_2_pt_V => fifo_out(7*NFIFOS+2).pt,
                     fifo_out_7_3_pt_V => fifo_out(7*NFIFOS+3).pt,
                     fifo_out_7_4_pt_V => fifo_out(7*NFIFOS+4).pt,
                     fifo_out_7_5_pt_V => fifo_out(7*NFIFOS+5).pt,
                     fifo_out_7_0_eta_V => fifo_out(7*NFIFOS+0).eta,
                     fifo_out_7_1_eta_V => fifo_out(7*NFIFOS+1).eta,
                     fifo_out_7_2_eta_V => fifo_out(7*NFIFOS+2).eta,
                     fifo_out_7_3_eta_V => fifo_out(7*NFIFOS+3).eta,
                     fifo_out_7_4_eta_V => fifo_out(7*NFIFOS+4).eta,
                     fifo_out_7_5_eta_V => fifo_out(7*NFIFOS+5).eta,
                     fifo_out_7_0_phi_V => fifo_out(7*NFIFOS+0).phi,
                     fifo_out_7_1_phi_V => fifo_out(7*NFIFOS+1).phi,
                     fifo_out_7_2_phi_V => fifo_out(7*NFIFOS+2).phi,
                     fifo_out_7_3_phi_V => fifo_out(7*NFIFOS+3).phi,
                     fifo_out_7_4_phi_V => fifo_out(7*NFIFOS+4).phi,
                     fifo_out_7_5_phi_V => fifo_out(7*NFIFOS+5).phi,
                     fifo_out_7_0_rest_V => fifo_out(7*NFIFOS+0).rest,
                     fifo_out_7_1_rest_V => fifo_out(7*NFIFOS+1).rest,
                     fifo_out_7_2_rest_V => fifo_out(7*NFIFOS+2).rest,
                     fifo_out_7_3_rest_V => fifo_out(7*NFIFOS+3).rest,
                     fifo_out_7_4_rest_V => fifo_out(7*NFIFOS+4).rest,
                     fifo_out_7_5_rest_V => fifo_out(7*NFIFOS+5).rest,
                     fifo_out_8_0_pt_V => fifo_out(8*NFIFOS+0).pt,
                     fifo_out_8_1_pt_V => fifo_out(8*NFIFOS+1).pt,
                     fifo_out_8_2_pt_V => fifo_out(8*NFIFOS+2).pt,
                     fifo_out_8_3_pt_V => fifo_out(8*NFIFOS+3).pt,
                     fifo_out_8_4_pt_V => fifo_out(8*NFIFOS+4).pt,
                     fifo_out_8_5_pt_V => fifo_out(8*NFIFOS+5).pt,
                     fifo_out_8_0_eta_V => fifo_out(8*NFIFOS+0).eta,
                     fifo_out_8_1_eta_V => fifo_out(8*NFIFOS+1).eta,
                     fifo_out_8_2_eta_V => fifo_out(8*NFIFOS+2).eta,
                     fifo_out_8_3_eta_V => fifo_out(8*NFIFOS+3).eta,
                     fifo_out_8_4_eta_V => fifo_out(8*NFIFOS+4).eta,
                     fifo_out_8_5_eta_V => fifo_out(8*NFIFOS+5).eta,
                     fifo_out_8_0_phi_V => fifo_out(8*NFIFOS+0).phi,
                     fifo_out_8_1_phi_V => fifo_out(8*NFIFOS+1).phi,
                     fifo_out_8_2_phi_V => fifo_out(8*NFIFOS+2).phi,
                     fifo_out_8_3_phi_V => fifo_out(8*NFIFOS+3).phi,
                     fifo_out_8_4_phi_V => fifo_out(8*NFIFOS+4).phi,
                     fifo_out_8_5_phi_V => fifo_out(8*NFIFOS+5).phi,
                     fifo_out_8_0_rest_V => fifo_out(8*NFIFOS+0).rest,
                     fifo_out_8_1_rest_V => fifo_out(8*NFIFOS+1).rest,
                     fifo_out_8_2_rest_V => fifo_out(8*NFIFOS+2).rest,
                     fifo_out_8_3_rest_V => fifo_out(8*NFIFOS+3).rest,
                     fifo_out_8_4_rest_V => fifo_out(8*NFIFOS+4).rest,
                     fifo_out_8_5_rest_V => fifo_out(8*NFIFOS+5).rest,
                     fifo_out_valid_0_0 => fifo_out_valid(0*NFIFOS+0),
                     fifo_out_valid_0_1 => fifo_out_valid(0*NFIFOS+1),
                     fifo_out_valid_0_2 => fifo_out_valid(0*NFIFOS+2),
                     fifo_out_valid_0_3 => fifo_out_valid(0*NFIFOS+3),
                     fifo_out_valid_0_4 => fifo_out_valid(0*NFIFOS+4),
                     fifo_out_valid_0_5 => fifo_out_valid(0*NFIFOS+5),
                     fifo_out_valid_1_0 => fifo_out_valid(1*NFIFOS+0),
                     fifo_out_valid_1_1 => fifo_out_valid(1*NFIFOS+1),
                     fifo_out_valid_1_2 => fifo_out_valid(1*NFIFOS+2),
                     fifo_out_valid_1_3 => fifo_out_valid(1*NFIFOS+3),
                     fifo_out_valid_1_4 => fifo_out_valid(1*NFIFOS+4),
                     fifo_out_valid_1_5 => fifo_out_valid(1*NFIFOS+5),
                     fifo_out_valid_2_0 => fifo_out_valid(2*NFIFOS+0),
                     fifo_out_valid_2_1 => fifo_out_valid(2*NFIFOS+1),
                     fifo_out_valid_2_2 => fifo_out_valid(2*NFIFOS+2),
                     fifo_out_valid_2_3 => fifo_out_valid(2*NFIFOS+3),
                     fifo_out_valid_2_4 => fifo_out_valid(2*NFIFOS+4),
                     fifo_out_valid_2_5 => fifo_out_valid(2*NFIFOS+5),
                     fifo_out_valid_3_0 => fifo_out_valid(3*NFIFOS+0),
                     fifo_out_valid_3_1 => fifo_out_valid(3*NFIFOS+1),
                     fifo_out_valid_3_2 => fifo_out_valid(3*NFIFOS+2),
                     fifo_out_valid_3_3 => fifo_out_valid(3*NFIFOS+3),
                     fifo_out_valid_3_4 => fifo_out_valid(3*NFIFOS+4),
                     fifo_out_valid_3_5 => fifo_out_valid(3*NFIFOS+5),
                     fifo_out_valid_4_0 => fifo_out_valid(4*NFIFOS+0),
                     fifo_out_valid_4_1 => fifo_out_valid(4*NFIFOS+1),
                     fifo_out_valid_4_2 => fifo_out_valid(4*NFIFOS+2),
                     fifo_out_valid_4_3 => fifo_out_valid(4*NFIFOS+3),
                     fifo_out_valid_4_4 => fifo_out_valid(4*NFIFOS+4),
                     fifo_out_valid_4_5 => fifo_out_valid(4*NFIFOS+5),
                     fifo_out_valid_5_0 => fifo_out_valid(5*NFIFOS+0),
                     fifo_out_valid_5_1 => fifo_out_valid(5*NFIFOS+1),
                     fifo_out_valid_5_2 => fifo_out_valid(5*NFIFOS+2),
                     fifo_out_valid_5_3 => fifo_out_valid(5*NFIFOS+3),
                     fifo_out_valid_5_4 => fifo_out_valid(5*NFIFOS+4),
                     fifo_out_valid_5_5 => fifo_out_valid(5*NFIFOS+5),
                     fifo_out_valid_6_0 => fifo_out_valid(6*NFIFOS+0),
                     fifo_out_valid_6_1 => fifo_out_valid(6*NFIFOS+1),
                     fifo_out_valid_6_2 => fifo_out_valid(6*NFIFOS+2),
                     fifo_out_valid_6_3 => fifo_out_valid(6*NFIFOS+3),
                     fifo_out_valid_6_4 => fifo_out_valid(6*NFIFOS+4),
                     fifo_out_valid_6_5 => fifo_out_valid(6*NFIFOS+5),
                     fifo_out_valid_7_0 => fifo_out_valid(7*NFIFOS+0),
                     fifo_out_valid_7_1 => fifo_out_valid(7*NFIFOS+1),
                     fifo_out_valid_7_2 => fifo_out_valid(7*NFIFOS+2),
                     fifo_out_valid_7_3 => fifo_out_valid(7*NFIFOS+3),
                     fifo_out_valid_7_4 => fifo_out_valid(7*NFIFOS+4),
                     fifo_out_valid_7_5 => fifo_out_valid(7*NFIFOS+5),
                     fifo_out_valid_8_0 => fifo_out_valid(8*NFIFOS+0),
                     fifo_out_valid_8_1 => fifo_out_valid(8*NFIFOS+1),
                     fifo_out_valid_8_2 => fifo_out_valid(8*NFIFOS+2),
                     fifo_out_valid_8_3 => fifo_out_valid(8*NFIFOS+3),
                     fifo_out_valid_8_4 => fifo_out_valid(8*NFIFOS+4),
                     fifo_out_valid_8_5 => fifo_out_valid(8*NFIFOS+5),
                     fifo_out_roll_0_0 => fifo_out_roll(0*NFIFOS+0),
                     fifo_out_roll_0_1 => fifo_out_roll(0*NFIFOS+1),
                     fifo_out_roll_0_2 => fifo_out_roll(0*NFIFOS+2),
                     fifo_out_roll_0_3 => fifo_out_roll(0*NFIFOS+3),
                     fifo_out_roll_0_4 => fifo_out_roll(0*NFIFOS+4),
                     fifo_out_roll_0_5 => fifo_out_roll(0*NFIFOS+5),
                     fifo_out_roll_1_0 => fifo_out_roll(1*NFIFOS+0),
                     fifo_out_roll_1_1 => fifo_out_roll(1*NFIFOS+1),
                     fifo_out_roll_1_2 => fifo_out_roll(1*NFIFOS+2),
                     fifo_out_roll_1_3 => fifo_out_roll(1*NFIFOS+3),
                     fifo_out_roll_1_4 => fifo_out_roll(1*NFIFOS+4),
                     fifo_out_roll_1_5 => fifo_out_roll(1*NFIFOS+5),
                     fifo_out_roll_2_0 => fifo_out_roll(2*NFIFOS+0),
                     fifo_out_roll_2_1 => fifo_out_roll(2*NFIFOS+1),
                     fifo_out_roll_2_2 => fifo_out_roll(2*NFIFOS+2),
                     fifo_out_roll_2_3 => fifo_out_roll(2*NFIFOS+3),
                     fifo_out_roll_2_4 => fifo_out_roll(2*NFIFOS+4),
                     fifo_out_roll_2_5 => fifo_out_roll(2*NFIFOS+5),
                     fifo_out_roll_3_0 => fifo_out_roll(3*NFIFOS+0),
                     fifo_out_roll_3_1 => fifo_out_roll(3*NFIFOS+1),
                     fifo_out_roll_3_2 => fifo_out_roll(3*NFIFOS+2),
                     fifo_out_roll_3_3 => fifo_out_roll(3*NFIFOS+3),
                     fifo_out_roll_3_4 => fifo_out_roll(3*NFIFOS+4),
                     fifo_out_roll_3_5 => fifo_out_roll(3*NFIFOS+5),
                     fifo_out_roll_4_0 => fifo_out_roll(4*NFIFOS+0),
                     fifo_out_roll_4_1 => fifo_out_roll(4*NFIFOS+1),
                     fifo_out_roll_4_2 => fifo_out_roll(4*NFIFOS+2),
                     fifo_out_roll_4_3 => fifo_out_roll(4*NFIFOS+3),
                     fifo_out_roll_4_4 => fifo_out_roll(4*NFIFOS+4),
                     fifo_out_roll_4_5 => fifo_out_roll(4*NFIFOS+5),
                     fifo_out_roll_5_0 => fifo_out_roll(5*NFIFOS+0),
                     fifo_out_roll_5_1 => fifo_out_roll(5*NFIFOS+1),
                     fifo_out_roll_5_2 => fifo_out_roll(5*NFIFOS+2),
                     fifo_out_roll_5_3 => fifo_out_roll(5*NFIFOS+3),
                     fifo_out_roll_5_4 => fifo_out_roll(5*NFIFOS+4),
                     fifo_out_roll_5_5 => fifo_out_roll(5*NFIFOS+5),
                     fifo_out_roll_6_0 => fifo_out_roll(6*NFIFOS+0),
                     fifo_out_roll_6_1 => fifo_out_roll(6*NFIFOS+1),
                     fifo_out_roll_6_2 => fifo_out_roll(6*NFIFOS+2),
                     fifo_out_roll_6_3 => fifo_out_roll(6*NFIFOS+3),
                     fifo_out_roll_6_4 => fifo_out_roll(6*NFIFOS+4),
                     fifo_out_roll_6_5 => fifo_out_roll(6*NFIFOS+5),
                     fifo_out_roll_7_0 => fifo_out_roll(7*NFIFOS+0),
                     fifo_out_roll_7_1 => fifo_out_roll(7*NFIFOS+1),
                     fifo_out_roll_7_2 => fifo_out_roll(7*NFIFOS+2),
                     fifo_out_roll_7_3 => fifo_out_roll(7*NFIFOS+3),
                     fifo_out_roll_7_4 => fifo_out_roll(7*NFIFOS+4),
                     fifo_out_roll_7_5 => fifo_out_roll(7*NFIFOS+5),
                     fifo_out_roll_8_0 => fifo_out_roll(8*NFIFOS+0),
                     fifo_out_roll_8_1 => fifo_out_roll(8*NFIFOS+1),
                     fifo_out_roll_8_2 => fifo_out_roll(8*NFIFOS+2),
                     fifo_out_roll_8_3 => fifo_out_roll(8*NFIFOS+3),
                     fifo_out_roll_8_4 => fifo_out_roll(8*NFIFOS+4),
                     fifo_out_roll_8_5 => fifo_out_roll(8*NFIFOS+5),
                     fifo_full_0_0 => fifo_out_full(0*NFIFOS+0),
                     fifo_full_0_1 => fifo_out_full(0*NFIFOS+1),
                     fifo_full_0_2 => fifo_out_full(0*NFIFOS+2),
                     fifo_full_0_3 => fifo_out_full(0*NFIFOS+3),
                     fifo_full_0_4 => fifo_out_full(0*NFIFOS+4),
                     fifo_full_0_5 => fifo_out_full(0*NFIFOS+5),
                     fifo_full_1_0 => fifo_out_full(1*NFIFOS+0),
                     fifo_full_1_1 => fifo_out_full(1*NFIFOS+1),
                     fifo_full_1_2 => fifo_out_full(1*NFIFOS+2),
                     fifo_full_1_3 => fifo_out_full(1*NFIFOS+3),
                     fifo_full_1_4 => fifo_out_full(1*NFIFOS+4),
                     fifo_full_1_5 => fifo_out_full(1*NFIFOS+5),
                     fifo_full_2_0 => fifo_out_full(2*NFIFOS+0),
                     fifo_full_2_1 => fifo_out_full(2*NFIFOS+1),
                     fifo_full_2_2 => fifo_out_full(2*NFIFOS+2),
                     fifo_full_2_3 => fifo_out_full(2*NFIFOS+3),
                     fifo_full_2_4 => fifo_out_full(2*NFIFOS+4),
                     fifo_full_2_5 => fifo_out_full(2*NFIFOS+5),
                     fifo_full_3_0 => fifo_out_full(3*NFIFOS+0),
                     fifo_full_3_1 => fifo_out_full(3*NFIFOS+1),
                     fifo_full_3_2 => fifo_out_full(3*NFIFOS+2),
                     fifo_full_3_3 => fifo_out_full(3*NFIFOS+3),
                     fifo_full_3_4 => fifo_out_full(3*NFIFOS+4),
                     fifo_full_3_5 => fifo_out_full(3*NFIFOS+5),
                     fifo_full_4_0 => fifo_out_full(4*NFIFOS+0),
                     fifo_full_4_1 => fifo_out_full(4*NFIFOS+1),
                     fifo_full_4_2 => fifo_out_full(4*NFIFOS+2),
                     fifo_full_4_3 => fifo_out_full(4*NFIFOS+3),
                     fifo_full_4_4 => fifo_out_full(4*NFIFOS+4),
                     fifo_full_4_5 => fifo_out_full(4*NFIFOS+5),
                     fifo_full_5_0 => fifo_out_full(5*NFIFOS+0),
                     fifo_full_5_1 => fifo_out_full(5*NFIFOS+1),
                     fifo_full_5_2 => fifo_out_full(5*NFIFOS+2),
                     fifo_full_5_3 => fifo_out_full(5*NFIFOS+3),
                     fifo_full_5_4 => fifo_out_full(5*NFIFOS+4),
                     fifo_full_5_5 => fifo_out_full(5*NFIFOS+5),
                     fifo_full_6_0 => fifo_out_full(6*NFIFOS+0),
                     fifo_full_6_1 => fifo_out_full(6*NFIFOS+1),
                     fifo_full_6_2 => fifo_out_full(6*NFIFOS+2),
                     fifo_full_6_3 => fifo_out_full(6*NFIFOS+3),
                     fifo_full_6_4 => fifo_out_full(6*NFIFOS+4),
                     fifo_full_6_5 => fifo_out_full(6*NFIFOS+5),
                     fifo_full_7_0 => fifo_out_full(7*NFIFOS+0),
                     fifo_full_7_1 => fifo_out_full(7*NFIFOS+1),
                     fifo_full_7_2 => fifo_out_full(7*NFIFOS+2),
                     fifo_full_7_3 => fifo_out_full(7*NFIFOS+3),
                     fifo_full_7_4 => fifo_out_full(7*NFIFOS+4),
                     fifo_full_7_5 => fifo_out_full(7*NFIFOS+5),
                     fifo_full_8_0 => fifo_out_full(8*NFIFOS+0),
                     fifo_full_8_1 => fifo_out_full(8*NFIFOS+1),
                     fifo_full_8_2 => fifo_out_full(8*NFIFOS+2),
                     fifo_full_8_3 => fifo_out_full(8*NFIFOS+3),
                     fifo_full_8_4 => fifo_out_full(8*NFIFOS+4),
                     fifo_full_8_5 => fifo_out_full(8*NFIFOS+5),
                     merged_out_0_0_pt_V => merged2_out(0*NFIFOS/2+0).pt,
                     merged_out_0_1_pt_V => merged2_out(0*NFIFOS/2+1).pt,
                     merged_out_0_2_pt_V => merged2_out(0*NFIFOS/2+2).pt,
                     merged_out_0_0_eta_V => merged2_out(0*NFIFOS/2+0).eta,
                     merged_out_0_1_eta_V => merged2_out(0*NFIFOS/2+1).eta,
                     merged_out_0_2_eta_V => merged2_out(0*NFIFOS/2+2).eta,
                     merged_out_0_0_phi_V => merged2_out(0*NFIFOS/2+0).phi,
                     merged_out_0_1_phi_V => merged2_out(0*NFIFOS/2+1).phi,
                     merged_out_0_2_phi_V => merged2_out(0*NFIFOS/2+2).phi,
                     merged_out_0_0_rest_V => merged2_out(0*NFIFOS/2+0).rest,
                     merged_out_0_1_rest_V => merged2_out(0*NFIFOS/2+1).rest,
                     merged_out_0_2_rest_V => merged2_out(0*NFIFOS/2+2).rest,
                     merged_out_1_0_pt_V => merged2_out(1*NFIFOS/2+0).pt,
                     merged_out_1_1_pt_V => merged2_out(1*NFIFOS/2+1).pt,
                     merged_out_1_2_pt_V => merged2_out(1*NFIFOS/2+2).pt,
                     merged_out_1_0_eta_V => merged2_out(1*NFIFOS/2+0).eta,
                     merged_out_1_1_eta_V => merged2_out(1*NFIFOS/2+1).eta,
                     merged_out_1_2_eta_V => merged2_out(1*NFIFOS/2+2).eta,
                     merged_out_1_0_phi_V => merged2_out(1*NFIFOS/2+0).phi,
                     merged_out_1_1_phi_V => merged2_out(1*NFIFOS/2+1).phi,
                     merged_out_1_2_phi_V => merged2_out(1*NFIFOS/2+2).phi,
                     merged_out_1_0_rest_V => merged2_out(1*NFIFOS/2+0).rest,
                     merged_out_1_1_rest_V => merged2_out(1*NFIFOS/2+1).rest,
                     merged_out_1_2_rest_V => merged2_out(1*NFIFOS/2+2).rest,
                     merged_out_2_0_pt_V => merged2_out(2*NFIFOS/2+0).pt,
                     merged_out_2_1_pt_V => merged2_out(2*NFIFOS/2+1).pt,
                     merged_out_2_2_pt_V => merged2_out(2*NFIFOS/2+2).pt,
                     merged_out_2_0_eta_V => merged2_out(2*NFIFOS/2+0).eta,
                     merged_out_2_1_eta_V => merged2_out(2*NFIFOS/2+1).eta,
                     merged_out_2_2_eta_V => merged2_out(2*NFIFOS/2+2).eta,
                     merged_out_2_0_phi_V => merged2_out(2*NFIFOS/2+0).phi,
                     merged_out_2_1_phi_V => merged2_out(2*NFIFOS/2+1).phi,
                     merged_out_2_2_phi_V => merged2_out(2*NFIFOS/2+2).phi,
                     merged_out_2_0_rest_V => merged2_out(2*NFIFOS/2+0).rest,
                     merged_out_2_1_rest_V => merged2_out(2*NFIFOS/2+1).rest,
                     merged_out_2_2_rest_V => merged2_out(2*NFIFOS/2+2).rest,
                     merged_out_3_0_pt_V => merged2_out(3*NFIFOS/2+0).pt,
                     merged_out_3_1_pt_V => merged2_out(3*NFIFOS/2+1).pt,
                     merged_out_3_2_pt_V => merged2_out(3*NFIFOS/2+2).pt,
                     merged_out_3_0_eta_V => merged2_out(3*NFIFOS/2+0).eta,
                     merged_out_3_1_eta_V => merged2_out(3*NFIFOS/2+1).eta,
                     merged_out_3_2_eta_V => merged2_out(3*NFIFOS/2+2).eta,
                     merged_out_3_0_phi_V => merged2_out(3*NFIFOS/2+0).phi,
                     merged_out_3_1_phi_V => merged2_out(3*NFIFOS/2+1).phi,
                     merged_out_3_2_phi_V => merged2_out(3*NFIFOS/2+2).phi,
                     merged_out_3_0_rest_V => merged2_out(3*NFIFOS/2+0).rest,
                     merged_out_3_1_rest_V => merged2_out(3*NFIFOS/2+1).rest,
                     merged_out_3_2_rest_V => merged2_out(3*NFIFOS/2+2).rest,
                     merged_out_4_0_pt_V => merged2_out(4*NFIFOS/2+0).pt,
                     merged_out_4_1_pt_V => merged2_out(4*NFIFOS/2+1).pt,
                     merged_out_4_2_pt_V => merged2_out(4*NFIFOS/2+2).pt,
                     merged_out_4_0_eta_V => merged2_out(4*NFIFOS/2+0).eta,
                     merged_out_4_1_eta_V => merged2_out(4*NFIFOS/2+1).eta,
                     merged_out_4_2_eta_V => merged2_out(4*NFIFOS/2+2).eta,
                     merged_out_4_0_phi_V => merged2_out(4*NFIFOS/2+0).phi,
                     merged_out_4_1_phi_V => merged2_out(4*NFIFOS/2+1).phi,
                     merged_out_4_2_phi_V => merged2_out(4*NFIFOS/2+2).phi,
                     merged_out_4_0_rest_V => merged2_out(4*NFIFOS/2+0).rest,
                     merged_out_4_1_rest_V => merged2_out(4*NFIFOS/2+1).rest,
                     merged_out_4_2_rest_V => merged2_out(4*NFIFOS/2+2).rest,
                     merged_out_5_0_pt_V => merged2_out(5*NFIFOS/2+0).pt,
                     merged_out_5_1_pt_V => merged2_out(5*NFIFOS/2+1).pt,
                     merged_out_5_2_pt_V => merged2_out(5*NFIFOS/2+2).pt,
                     merged_out_5_0_eta_V => merged2_out(5*NFIFOS/2+0).eta,
                     merged_out_5_1_eta_V => merged2_out(5*NFIFOS/2+1).eta,
                     merged_out_5_2_eta_V => merged2_out(5*NFIFOS/2+2).eta,
                     merged_out_5_0_phi_V => merged2_out(5*NFIFOS/2+0).phi,
                     merged_out_5_1_phi_V => merged2_out(5*NFIFOS/2+1).phi,
                     merged_out_5_2_phi_V => merged2_out(5*NFIFOS/2+2).phi,
                     merged_out_5_0_rest_V => merged2_out(5*NFIFOS/2+0).rest,
                     merged_out_5_1_rest_V => merged2_out(5*NFIFOS/2+1).rest,
                     merged_out_5_2_rest_V => merged2_out(5*NFIFOS/2+2).rest,
                     merged_out_6_0_pt_V => merged2_out(6*NFIFOS/2+0).pt,
                     merged_out_6_1_pt_V => merged2_out(6*NFIFOS/2+1).pt,
                     merged_out_6_2_pt_V => merged2_out(6*NFIFOS/2+2).pt,
                     merged_out_6_0_eta_V => merged2_out(6*NFIFOS/2+0).eta,
                     merged_out_6_1_eta_V => merged2_out(6*NFIFOS/2+1).eta,
                     merged_out_6_2_eta_V => merged2_out(6*NFIFOS/2+2).eta,
                     merged_out_6_0_phi_V => merged2_out(6*NFIFOS/2+0).phi,
                     merged_out_6_1_phi_V => merged2_out(6*NFIFOS/2+1).phi,
                     merged_out_6_2_phi_V => merged2_out(6*NFIFOS/2+2).phi,
                     merged_out_6_0_rest_V => merged2_out(6*NFIFOS/2+0).rest,
                     merged_out_6_1_rest_V => merged2_out(6*NFIFOS/2+1).rest,
                     merged_out_6_2_rest_V => merged2_out(6*NFIFOS/2+2).rest,
                     merged_out_7_0_pt_V => merged2_out(7*NFIFOS/2+0).pt,
                     merged_out_7_1_pt_V => merged2_out(7*NFIFOS/2+1).pt,
                     merged_out_7_2_pt_V => merged2_out(7*NFIFOS/2+2).pt,
                     merged_out_7_0_eta_V => merged2_out(7*NFIFOS/2+0).eta,
                     merged_out_7_1_eta_V => merged2_out(7*NFIFOS/2+1).eta,
                     merged_out_7_2_eta_V => merged2_out(7*NFIFOS/2+2).eta,
                     merged_out_7_0_phi_V => merged2_out(7*NFIFOS/2+0).phi,
                     merged_out_7_1_phi_V => merged2_out(7*NFIFOS/2+1).phi,
                     merged_out_7_2_phi_V => merged2_out(7*NFIFOS/2+2).phi,
                     merged_out_7_0_rest_V => merged2_out(7*NFIFOS/2+0).rest,
                     merged_out_7_1_rest_V => merged2_out(7*NFIFOS/2+1).rest,
                     merged_out_7_2_rest_V => merged2_out(7*NFIFOS/2+2).rest,
                     merged_out_8_0_pt_V => merged2_out(8*NFIFOS/2+0).pt,
                     merged_out_8_1_pt_V => merged2_out(8*NFIFOS/2+1).pt,
                     merged_out_8_2_pt_V => merged2_out(8*NFIFOS/2+2).pt,
                     merged_out_8_0_eta_V => merged2_out(8*NFIFOS/2+0).eta,
                     merged_out_8_1_eta_V => merged2_out(8*NFIFOS/2+1).eta,
                     merged_out_8_2_eta_V => merged2_out(8*NFIFOS/2+2).eta,
                     merged_out_8_0_phi_V => merged2_out(8*NFIFOS/2+0).phi,
                     merged_out_8_1_phi_V => merged2_out(8*NFIFOS/2+1).phi,
                     merged_out_8_2_phi_V => merged2_out(8*NFIFOS/2+2).phi,
                     merged_out_8_0_rest_V => merged2_out(8*NFIFOS/2+0).rest,
                     merged_out_8_1_rest_V => merged2_out(8*NFIFOS/2+1).rest,
                     merged_out_8_2_rest_V => merged2_out(8*NFIFOS/2+2).rest,
                     merged_out_valid_0_0 => merged2_out_valid(0*NFIFOS/2+0),
                     merged_out_valid_0_1 => merged2_out_valid(0*NFIFOS/2+1),
                     merged_out_valid_0_2 => merged2_out_valid(0*NFIFOS/2+2),
                     merged_out_valid_1_0 => merged2_out_valid(1*NFIFOS/2+0),
                     merged_out_valid_1_1 => merged2_out_valid(1*NFIFOS/2+1),
                     merged_out_valid_1_2 => merged2_out_valid(1*NFIFOS/2+2),
                     merged_out_valid_2_0 => merged2_out_valid(2*NFIFOS/2+0),
                     merged_out_valid_2_1 => merged2_out_valid(2*NFIFOS/2+1),
                     merged_out_valid_2_2 => merged2_out_valid(2*NFIFOS/2+2),
                     merged_out_valid_3_0 => merged2_out_valid(3*NFIFOS/2+0),
                     merged_out_valid_3_1 => merged2_out_valid(3*NFIFOS/2+1),
                     merged_out_valid_3_2 => merged2_out_valid(3*NFIFOS/2+2),
                     merged_out_valid_4_0 => merged2_out_valid(4*NFIFOS/2+0),
                     merged_out_valid_4_1 => merged2_out_valid(4*NFIFOS/2+1),
                     merged_out_valid_4_2 => merged2_out_valid(4*NFIFOS/2+2),
                     merged_out_valid_5_0 => merged2_out_valid(5*NFIFOS/2+0),
                     merged_out_valid_5_1 => merged2_out_valid(5*NFIFOS/2+1),
                     merged_out_valid_5_2 => merged2_out_valid(5*NFIFOS/2+2),
                     merged_out_valid_6_0 => merged2_out_valid(6*NFIFOS/2+0),
                     merged_out_valid_6_1 => merged2_out_valid(6*NFIFOS/2+1),
                     merged_out_valid_6_2 => merged2_out_valid(6*NFIFOS/2+2),
                     merged_out_valid_7_0 => merged2_out_valid(7*NFIFOS/2+0),
                     merged_out_valid_7_1 => merged2_out_valid(7*NFIFOS/2+1),
                     merged_out_valid_7_2 => merged2_out_valid(7*NFIFOS/2+2),
                     merged_out_valid_8_0 => merged2_out_valid(8*NFIFOS/2+0),
                     merged_out_valid_8_1 => merged2_out_valid(8*NFIFOS/2+1),
                     merged_out_valid_8_2 => merged2_out_valid(8*NFIFOS/2+2),
                     merged_out_roll_0_0 => merged2_out_roll(0*NFIFOS/2+0),
                     merged_out_roll_0_1 => merged2_out_roll(0*NFIFOS/2+1),
                     merged_out_roll_0_2 => merged2_out_roll(0*NFIFOS/2+2),
                     merged_out_roll_1_0 => merged2_out_roll(1*NFIFOS/2+0),
                     merged_out_roll_1_1 => merged2_out_roll(1*NFIFOS/2+1),
                     merged_out_roll_1_2 => merged2_out_roll(1*NFIFOS/2+2),
                     merged_out_roll_2_0 => merged2_out_roll(2*NFIFOS/2+0),
                     merged_out_roll_2_1 => merged2_out_roll(2*NFIFOS/2+1),
                     merged_out_roll_2_2 => merged2_out_roll(2*NFIFOS/2+2),
                     merged_out_roll_3_0 => merged2_out_roll(3*NFIFOS/2+0),
                     merged_out_roll_3_1 => merged2_out_roll(3*NFIFOS/2+1),
                     merged_out_roll_3_2 => merged2_out_roll(3*NFIFOS/2+2),
                     merged_out_roll_4_0 => merged2_out_roll(4*NFIFOS/2+0),
                     merged_out_roll_4_1 => merged2_out_roll(4*NFIFOS/2+1),
                     merged_out_roll_4_2 => merged2_out_roll(4*NFIFOS/2+2),
                     merged_out_roll_5_0 => merged2_out_roll(5*NFIFOS/2+0),
                     merged_out_roll_5_1 => merged2_out_roll(5*NFIFOS/2+1),
                     merged_out_roll_5_2 => merged2_out_roll(5*NFIFOS/2+2),
                     merged_out_roll_6_0 => merged2_out_roll(6*NFIFOS/2+0),
                     merged_out_roll_6_1 => merged2_out_roll(6*NFIFOS/2+1),
                     merged_out_roll_6_2 => merged2_out_roll(6*NFIFOS/2+2),
                     merged_out_roll_7_0 => merged2_out_roll(7*NFIFOS/2+0),
                     merged_out_roll_7_1 => merged2_out_roll(7*NFIFOS/2+1),
                     merged_out_roll_7_2 => merged2_out_roll(7*NFIFOS/2+2),
                     merged_out_roll_8_0 => merged2_out_roll(8*NFIFOS/2+0),
                     merged_out_roll_8_1 => merged2_out_roll(8*NFIFOS/2+1),
                     merged_out_roll_8_2 => merged2_out_roll(8*NFIFOS/2+2),
                     merged_full_0_0 => merged2_full(0*NFIFOS/2+0),
                     merged_full_0_1 => merged2_full(0*NFIFOS/2+1),
                     merged_full_0_2 => merged2_full(0*NFIFOS/2+2),
                     merged_full_1_0 => merged2_full(1*NFIFOS/2+0),
                     merged_full_1_1 => merged2_full(1*NFIFOS/2+1),
                     merged_full_1_2 => merged2_full(1*NFIFOS/2+2),
                     merged_full_2_0 => merged2_full(2*NFIFOS/2+0),
                     merged_full_2_1 => merged2_full(2*NFIFOS/2+1),
                     merged_full_2_2 => merged2_full(2*NFIFOS/2+2),
                     merged_full_3_0 => merged2_full(3*NFIFOS/2+0),
                     merged_full_3_1 => merged2_full(3*NFIFOS/2+1),
                     merged_full_3_2 => merged2_full(3*NFIFOS/2+2),
                     merged_full_4_0 => merged2_full(4*NFIFOS/2+0),
                     merged_full_4_1 => merged2_full(4*NFIFOS/2+1),
                     merged_full_4_2 => merged2_full(4*NFIFOS/2+2),
                     merged_full_5_0 => merged2_full(5*NFIFOS/2+0),
                     merged_full_5_1 => merged2_full(5*NFIFOS/2+1),
                     merged_full_5_2 => merged2_full(5*NFIFOS/2+2),
                     merged_full_6_0 => merged2_full(6*NFIFOS/2+0),
                     merged_full_6_1 => merged2_full(6*NFIFOS/2+1),
                     merged_full_6_2 => merged2_full(6*NFIFOS/2+2),
                     merged_full_7_0 => merged2_full(7*NFIFOS/2+0),
                     merged_full_7_1 => merged2_full(7*NFIFOS/2+1),
                     merged_full_7_2 => merged2_full(7*NFIFOS/2+2),
                     merged_full_8_0 => merged2_full(8*NFIFOS/2+0),
                     merged_full_8_1 => merged2_full(8*NFIFOS/2+1),
                     merged_full_8_2 => merged2_full(8*NFIFOS/2+2)
                 );

    merge3_slice : entity work.router_merge3_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     merged_out_0_0_pt_V => merged2_out(0*NFIFOS/2+0).pt,
                     merged_out_0_1_pt_V => merged2_out(0*NFIFOS/2+1).pt,
                     merged_out_0_2_pt_V => merged2_out(0*NFIFOS/2+2).pt,
                     merged_out_0_0_eta_V => merged2_out(0*NFIFOS/2+0).eta,
                     merged_out_0_1_eta_V => merged2_out(0*NFIFOS/2+1).eta,
                     merged_out_0_2_eta_V => merged2_out(0*NFIFOS/2+2).eta,
                     merged_out_0_0_phi_V => merged2_out(0*NFIFOS/2+0).phi,
                     merged_out_0_1_phi_V => merged2_out(0*NFIFOS/2+1).phi,
                     merged_out_0_2_phi_V => merged2_out(0*NFIFOS/2+2).phi,
                     merged_out_0_0_rest_V => merged2_out(0*NFIFOS/2+0).rest,
                     merged_out_0_1_rest_V => merged2_out(0*NFIFOS/2+1).rest,
                     merged_out_0_2_rest_V => merged2_out(0*NFIFOS/2+2).rest,
                     merged_out_1_0_pt_V => merged2_out(1*NFIFOS/2+0).pt,
                     merged_out_1_1_pt_V => merged2_out(1*NFIFOS/2+1).pt,
                     merged_out_1_2_pt_V => merged2_out(1*NFIFOS/2+2).pt,
                     merged_out_1_0_eta_V => merged2_out(1*NFIFOS/2+0).eta,
                     merged_out_1_1_eta_V => merged2_out(1*NFIFOS/2+1).eta,
                     merged_out_1_2_eta_V => merged2_out(1*NFIFOS/2+2).eta,
                     merged_out_1_0_phi_V => merged2_out(1*NFIFOS/2+0).phi,
                     merged_out_1_1_phi_V => merged2_out(1*NFIFOS/2+1).phi,
                     merged_out_1_2_phi_V => merged2_out(1*NFIFOS/2+2).phi,
                     merged_out_1_0_rest_V => merged2_out(1*NFIFOS/2+0).rest,
                     merged_out_1_1_rest_V => merged2_out(1*NFIFOS/2+1).rest,
                     merged_out_1_2_rest_V => merged2_out(1*NFIFOS/2+2).rest,
                     merged_out_2_0_pt_V => merged2_out(2*NFIFOS/2+0).pt,
                     merged_out_2_1_pt_V => merged2_out(2*NFIFOS/2+1).pt,
                     merged_out_2_2_pt_V => merged2_out(2*NFIFOS/2+2).pt,
                     merged_out_2_0_eta_V => merged2_out(2*NFIFOS/2+0).eta,
                     merged_out_2_1_eta_V => merged2_out(2*NFIFOS/2+1).eta,
                     merged_out_2_2_eta_V => merged2_out(2*NFIFOS/2+2).eta,
                     merged_out_2_0_phi_V => merged2_out(2*NFIFOS/2+0).phi,
                     merged_out_2_1_phi_V => merged2_out(2*NFIFOS/2+1).phi,
                     merged_out_2_2_phi_V => merged2_out(2*NFIFOS/2+2).phi,
                     merged_out_2_0_rest_V => merged2_out(2*NFIFOS/2+0).rest,
                     merged_out_2_1_rest_V => merged2_out(2*NFIFOS/2+1).rest,
                     merged_out_2_2_rest_V => merged2_out(2*NFIFOS/2+2).rest,
                     merged_out_3_0_pt_V => merged2_out(3*NFIFOS/2+0).pt,
                     merged_out_3_1_pt_V => merged2_out(3*NFIFOS/2+1).pt,
                     merged_out_3_2_pt_V => merged2_out(3*NFIFOS/2+2).pt,
                     merged_out_3_0_eta_V => merged2_out(3*NFIFOS/2+0).eta,
                     merged_out_3_1_eta_V => merged2_out(3*NFIFOS/2+1).eta,
                     merged_out_3_2_eta_V => merged2_out(3*NFIFOS/2+2).eta,
                     merged_out_3_0_phi_V => merged2_out(3*NFIFOS/2+0).phi,
                     merged_out_3_1_phi_V => merged2_out(3*NFIFOS/2+1).phi,
                     merged_out_3_2_phi_V => merged2_out(3*NFIFOS/2+2).phi,
                     merged_out_3_0_rest_V => merged2_out(3*NFIFOS/2+0).rest,
                     merged_out_3_1_rest_V => merged2_out(3*NFIFOS/2+1).rest,
                     merged_out_3_2_rest_V => merged2_out(3*NFIFOS/2+2).rest,
                     merged_out_4_0_pt_V => merged2_out(4*NFIFOS/2+0).pt,
                     merged_out_4_1_pt_V => merged2_out(4*NFIFOS/2+1).pt,
                     merged_out_4_2_pt_V => merged2_out(4*NFIFOS/2+2).pt,
                     merged_out_4_0_eta_V => merged2_out(4*NFIFOS/2+0).eta,
                     merged_out_4_1_eta_V => merged2_out(4*NFIFOS/2+1).eta,
                     merged_out_4_2_eta_V => merged2_out(4*NFIFOS/2+2).eta,
                     merged_out_4_0_phi_V => merged2_out(4*NFIFOS/2+0).phi,
                     merged_out_4_1_phi_V => merged2_out(4*NFIFOS/2+1).phi,
                     merged_out_4_2_phi_V => merged2_out(4*NFIFOS/2+2).phi,
                     merged_out_4_0_rest_V => merged2_out(4*NFIFOS/2+0).rest,
                     merged_out_4_1_rest_V => merged2_out(4*NFIFOS/2+1).rest,
                     merged_out_4_2_rest_V => merged2_out(4*NFIFOS/2+2).rest,
                     merged_out_5_0_pt_V => merged2_out(5*NFIFOS/2+0).pt,
                     merged_out_5_1_pt_V => merged2_out(5*NFIFOS/2+1).pt,
                     merged_out_5_2_pt_V => merged2_out(5*NFIFOS/2+2).pt,
                     merged_out_5_0_eta_V => merged2_out(5*NFIFOS/2+0).eta,
                     merged_out_5_1_eta_V => merged2_out(5*NFIFOS/2+1).eta,
                     merged_out_5_2_eta_V => merged2_out(5*NFIFOS/2+2).eta,
                     merged_out_5_0_phi_V => merged2_out(5*NFIFOS/2+0).phi,
                     merged_out_5_1_phi_V => merged2_out(5*NFIFOS/2+1).phi,
                     merged_out_5_2_phi_V => merged2_out(5*NFIFOS/2+2).phi,
                     merged_out_5_0_rest_V => merged2_out(5*NFIFOS/2+0).rest,
                     merged_out_5_1_rest_V => merged2_out(5*NFIFOS/2+1).rest,
                     merged_out_5_2_rest_V => merged2_out(5*NFIFOS/2+2).rest,
                     merged_out_6_0_pt_V => merged2_out(6*NFIFOS/2+0).pt,
                     merged_out_6_1_pt_V => merged2_out(6*NFIFOS/2+1).pt,
                     merged_out_6_2_pt_V => merged2_out(6*NFIFOS/2+2).pt,
                     merged_out_6_0_eta_V => merged2_out(6*NFIFOS/2+0).eta,
                     merged_out_6_1_eta_V => merged2_out(6*NFIFOS/2+1).eta,
                     merged_out_6_2_eta_V => merged2_out(6*NFIFOS/2+2).eta,
                     merged_out_6_0_phi_V => merged2_out(6*NFIFOS/2+0).phi,
                     merged_out_6_1_phi_V => merged2_out(6*NFIFOS/2+1).phi,
                     merged_out_6_2_phi_V => merged2_out(6*NFIFOS/2+2).phi,
                     merged_out_6_0_rest_V => merged2_out(6*NFIFOS/2+0).rest,
                     merged_out_6_1_rest_V => merged2_out(6*NFIFOS/2+1).rest,
                     merged_out_6_2_rest_V => merged2_out(6*NFIFOS/2+2).rest,
                     merged_out_7_0_pt_V => merged2_out(7*NFIFOS/2+0).pt,
                     merged_out_7_1_pt_V => merged2_out(7*NFIFOS/2+1).pt,
                     merged_out_7_2_pt_V => merged2_out(7*NFIFOS/2+2).pt,
                     merged_out_7_0_eta_V => merged2_out(7*NFIFOS/2+0).eta,
                     merged_out_7_1_eta_V => merged2_out(7*NFIFOS/2+1).eta,
                     merged_out_7_2_eta_V => merged2_out(7*NFIFOS/2+2).eta,
                     merged_out_7_0_phi_V => merged2_out(7*NFIFOS/2+0).phi,
                     merged_out_7_1_phi_V => merged2_out(7*NFIFOS/2+1).phi,
                     merged_out_7_2_phi_V => merged2_out(7*NFIFOS/2+2).phi,
                     merged_out_7_0_rest_V => merged2_out(7*NFIFOS/2+0).rest,
                     merged_out_7_1_rest_V => merged2_out(7*NFIFOS/2+1).rest,
                     merged_out_7_2_rest_V => merged2_out(7*NFIFOS/2+2).rest,
                     merged_out_8_0_pt_V => merged2_out(8*NFIFOS/2+0).pt,
                     merged_out_8_1_pt_V => merged2_out(8*NFIFOS/2+1).pt,
                     merged_out_8_2_pt_V => merged2_out(8*NFIFOS/2+2).pt,
                     merged_out_8_0_eta_V => merged2_out(8*NFIFOS/2+0).eta,
                     merged_out_8_1_eta_V => merged2_out(8*NFIFOS/2+1).eta,
                     merged_out_8_2_eta_V => merged2_out(8*NFIFOS/2+2).eta,
                     merged_out_8_0_phi_V => merged2_out(8*NFIFOS/2+0).phi,
                     merged_out_8_1_phi_V => merged2_out(8*NFIFOS/2+1).phi,
                     merged_out_8_2_phi_V => merged2_out(8*NFIFOS/2+2).phi,
                     merged_out_8_0_rest_V => merged2_out(8*NFIFOS/2+0).rest,
                     merged_out_8_1_rest_V => merged2_out(8*NFIFOS/2+1).rest,
                     merged_out_8_2_rest_V => merged2_out(8*NFIFOS/2+2).rest,
                     merged_out_valid_0_0 => merged2_out_valid(0*NFIFOS/2+0),
                     merged_out_valid_0_1 => merged2_out_valid(0*NFIFOS/2+1),
                     merged_out_valid_0_2 => merged2_out_valid(0*NFIFOS/2+2),
                     merged_out_valid_1_0 => merged2_out_valid(1*NFIFOS/2+0),
                     merged_out_valid_1_1 => merged2_out_valid(1*NFIFOS/2+1),
                     merged_out_valid_1_2 => merged2_out_valid(1*NFIFOS/2+2),
                     merged_out_valid_2_0 => merged2_out_valid(2*NFIFOS/2+0),
                     merged_out_valid_2_1 => merged2_out_valid(2*NFIFOS/2+1),
                     merged_out_valid_2_2 => merged2_out_valid(2*NFIFOS/2+2),
                     merged_out_valid_3_0 => merged2_out_valid(3*NFIFOS/2+0),
                     merged_out_valid_3_1 => merged2_out_valid(3*NFIFOS/2+1),
                     merged_out_valid_3_2 => merged2_out_valid(3*NFIFOS/2+2),
                     merged_out_valid_4_0 => merged2_out_valid(4*NFIFOS/2+0),
                     merged_out_valid_4_1 => merged2_out_valid(4*NFIFOS/2+1),
                     merged_out_valid_4_2 => merged2_out_valid(4*NFIFOS/2+2),
                     merged_out_valid_5_0 => merged2_out_valid(5*NFIFOS/2+0),
                     merged_out_valid_5_1 => merged2_out_valid(5*NFIFOS/2+1),
                     merged_out_valid_5_2 => merged2_out_valid(5*NFIFOS/2+2),
                     merged_out_valid_6_0 => merged2_out_valid(6*NFIFOS/2+0),
                     merged_out_valid_6_1 => merged2_out_valid(6*NFIFOS/2+1),
                     merged_out_valid_6_2 => merged2_out_valid(6*NFIFOS/2+2),
                     merged_out_valid_7_0 => merged2_out_valid(7*NFIFOS/2+0),
                     merged_out_valid_7_1 => merged2_out_valid(7*NFIFOS/2+1),
                     merged_out_valid_7_2 => merged2_out_valid(7*NFIFOS/2+2),
                     merged_out_valid_8_0 => merged2_out_valid(8*NFIFOS/2+0),
                     merged_out_valid_8_1 => merged2_out_valid(8*NFIFOS/2+1),
                     merged_out_valid_8_2 => merged2_out_valid(8*NFIFOS/2+2),
                     merged_out_roll_0_0 => merged2_out_roll(0*NFIFOS/2+0),
                     merged_out_roll_0_1 => merged2_out_roll(0*NFIFOS/2+1),
                     merged_out_roll_0_2 => merged2_out_roll(0*NFIFOS/2+2),
                     merged_out_roll_1_0 => merged2_out_roll(1*NFIFOS/2+0),
                     merged_out_roll_1_1 => merged2_out_roll(1*NFIFOS/2+1),
                     merged_out_roll_1_2 => merged2_out_roll(1*NFIFOS/2+2),
                     merged_out_roll_2_0 => merged2_out_roll(2*NFIFOS/2+0),
                     merged_out_roll_2_1 => merged2_out_roll(2*NFIFOS/2+1),
                     merged_out_roll_2_2 => merged2_out_roll(2*NFIFOS/2+2),
                     merged_out_roll_3_0 => merged2_out_roll(3*NFIFOS/2+0),
                     merged_out_roll_3_1 => merged2_out_roll(3*NFIFOS/2+1),
                     merged_out_roll_3_2 => merged2_out_roll(3*NFIFOS/2+2),
                     merged_out_roll_4_0 => merged2_out_roll(4*NFIFOS/2+0),
                     merged_out_roll_4_1 => merged2_out_roll(4*NFIFOS/2+1),
                     merged_out_roll_4_2 => merged2_out_roll(4*NFIFOS/2+2),
                     merged_out_roll_5_0 => merged2_out_roll(5*NFIFOS/2+0),
                     merged_out_roll_5_1 => merged2_out_roll(5*NFIFOS/2+1),
                     merged_out_roll_5_2 => merged2_out_roll(5*NFIFOS/2+2),
                     merged_out_roll_6_0 => merged2_out_roll(6*NFIFOS/2+0),
                     merged_out_roll_6_1 => merged2_out_roll(6*NFIFOS/2+1),
                     merged_out_roll_6_2 => merged2_out_roll(6*NFIFOS/2+2),
                     merged_out_roll_7_0 => merged2_out_roll(7*NFIFOS/2+0),
                     merged_out_roll_7_1 => merged2_out_roll(7*NFIFOS/2+1),
                     merged_out_roll_7_2 => merged2_out_roll(7*NFIFOS/2+2),
                     merged_out_roll_8_0 => merged2_out_roll(8*NFIFOS/2+0),
                     merged_out_roll_8_1 => merged2_out_roll(8*NFIFOS/2+1),
                     merged_out_roll_8_2 => merged2_out_roll(8*NFIFOS/2+2),
                     merged_full_0_0 => merged2_full(0*NFIFOS/2+0),
                     merged_full_0_1 => merged2_full(0*NFIFOS/2+1),
                     merged_full_0_2 => merged2_full(0*NFIFOS/2+2),
                     merged_full_1_0 => merged2_full(1*NFIFOS/2+0),
                     merged_full_1_1 => merged2_full(1*NFIFOS/2+1),
                     merged_full_1_2 => merged2_full(1*NFIFOS/2+2),
                     merged_full_2_0 => merged2_full(2*NFIFOS/2+0),
                     merged_full_2_1 => merged2_full(2*NFIFOS/2+1),
                     merged_full_2_2 => merged2_full(2*NFIFOS/2+2),
                     merged_full_3_0 => merged2_full(3*NFIFOS/2+0),
                     merged_full_3_1 => merged2_full(3*NFIFOS/2+1),
                     merged_full_3_2 => merged2_full(3*NFIFOS/2+2),
                     merged_full_4_0 => merged2_full(4*NFIFOS/2+0),
                     merged_full_4_1 => merged2_full(4*NFIFOS/2+1),
                     merged_full_4_2 => merged2_full(4*NFIFOS/2+2),
                     merged_full_5_0 => merged2_full(5*NFIFOS/2+0),
                     merged_full_5_1 => merged2_full(5*NFIFOS/2+1),
                     merged_full_5_2 => merged2_full(5*NFIFOS/2+2),
                     merged_full_6_0 => merged2_full(6*NFIFOS/2+0),
                     merged_full_6_1 => merged2_full(6*NFIFOS/2+1),
                     merged_full_6_2 => merged2_full(6*NFIFOS/2+2),
                     merged_full_7_0 => merged2_full(7*NFIFOS/2+0),
                     merged_full_7_1 => merged2_full(7*NFIFOS/2+1),
                     merged_full_7_2 => merged2_full(7*NFIFOS/2+2),
                     merged_full_8_0 => merged2_full(8*NFIFOS/2+0),
                     merged_full_8_1 => merged2_full(8*NFIFOS/2+1),
                     merged_full_8_2 => merged2_full(8*NFIFOS/2+2),
                     merged3_out_0_pt_V => merged_out(0).pt,
                     merged3_out_0_eta_V => merged_out(0).eta,
                     merged3_out_0_phi_V => merged_out(0).phi,
                     merged3_out_0_rest_V => merged_out(0).rest,
                     merged3_out_1_pt_V => merged_out(1).pt,
                     merged3_out_1_eta_V => merged_out(1).eta,
                     merged3_out_1_phi_V => merged_out(1).phi,
                     merged3_out_1_rest_V => merged_out(1).rest,
                     merged3_out_2_pt_V => merged_out(2).pt,
                     merged3_out_2_eta_V => merged_out(2).eta,
                     merged3_out_2_phi_V => merged_out(2).phi,
                     merged3_out_2_rest_V => merged_out(2).rest,
                     merged3_out_3_pt_V => merged_out(3).pt,
                     merged3_out_3_eta_V => merged_out(3).eta,
                     merged3_out_3_phi_V => merged_out(3).phi,
                     merged3_out_3_rest_V => merged_out(3).rest,
                     merged3_out_4_pt_V => merged_out(4).pt,
                     merged3_out_4_eta_V => merged_out(4).eta,
                     merged3_out_4_phi_V => merged_out(4).phi,
                     merged3_out_4_rest_V => merged_out(4).rest,
                     merged3_out_5_pt_V => merged_out(5).pt,
                     merged3_out_5_eta_V => merged_out(5).eta,
                     merged3_out_5_phi_V => merged_out(5).phi,
                     merged3_out_5_rest_V => merged_out(5).rest,
                     merged3_out_6_pt_V => merged_out(6).pt,
                     merged3_out_6_eta_V => merged_out(6).eta,
                     merged3_out_6_phi_V => merged_out(6).phi,
                     merged3_out_6_rest_V => merged_out(6).rest,
                     merged3_out_7_pt_V => merged_out(7).pt,
                     merged3_out_7_eta_V => merged_out(7).eta,
                     merged3_out_7_phi_V => merged_out(7).phi,
                     merged3_out_7_rest_V => merged_out(7).rest,
                     merged3_out_8_pt_V => merged_out(8).pt,
                     merged3_out_8_eta_V => merged_out(8).eta,
                     merged3_out_8_phi_V => merged_out(8).phi,
                     merged3_out_8_rest_V => merged_out(8).rest,
                     merged3_out_valid_0 => merged_out_valid(0),
                     merged3_out_valid_1 => merged_out_valid(1),
                     merged3_out_valid_2 => merged_out_valid(2),
                     merged3_out_valid_3 => merged_out_valid(3),
                     merged3_out_valid_4 => merged_out_valid(4),
                     merged3_out_valid_5 => merged_out_valid(5),
                     merged3_out_valid_6 => merged_out_valid(6),
                     merged3_out_valid_7 => merged_out_valid(7),
                     merged3_out_valid_8 => merged_out_valid(8),
                     merged3_out_roll_0 => merged_out_roll(0),
                     merged3_out_roll_1 => merged_out_roll(1),
                     merged3_out_roll_2 => merged_out_roll(2),
                     merged3_out_roll_3 => merged_out_roll(3),
                     merged3_out_roll_4 => merged_out_roll(4),
                     merged3_out_roll_5 => merged_out_roll(5),
                     merged3_out_roll_6 => merged_out_roll(6),
                     merged3_out_roll_7 => merged_out_roll(7),
                     merged3_out_roll_8 => merged_out_roll(8)
                 );


    output_slice : entity work.router_full_output_slice
            port map(ap_clk => ap_clk, 
                     ap_rst => ap_rst,
                     ap_start => '1',
                     ap_done => open,
                     ap_ready => open,
                     merged3_out_0_pt_V => merged_out(0).pt,
                     merged3_out_0_eta_V => merged_out(0).eta,
                     merged3_out_0_phi_V => merged_out(0).phi,
                     merged3_out_0_rest_V => merged_out(0).rest,
                     merged3_out_1_pt_V => merged_out(1).pt,
                     merged3_out_1_eta_V => merged_out(1).eta,
                     merged3_out_1_phi_V => merged_out(1).phi,
                     merged3_out_1_rest_V => merged_out(1).rest,
                     merged3_out_2_pt_V => merged_out(2).pt,
                     merged3_out_2_eta_V => merged_out(2).eta,
                     merged3_out_2_phi_V => merged_out(2).phi,
                     merged3_out_2_rest_V => merged_out(2).rest,
                     merged3_out_3_pt_V => merged_out(3).pt,
                     merged3_out_3_eta_V => merged_out(3).eta,
                     merged3_out_3_phi_V => merged_out(3).phi,
                     merged3_out_3_rest_V => merged_out(3).rest,
                     merged3_out_4_pt_V => merged_out(4).pt,
                     merged3_out_4_eta_V => merged_out(4).eta,
                     merged3_out_4_phi_V => merged_out(4).phi,
                     merged3_out_4_rest_V => merged_out(4).rest,
                     merged3_out_5_pt_V => merged_out(5).pt,
                     merged3_out_5_eta_V => merged_out(5).eta,
                     merged3_out_5_phi_V => merged_out(5).phi,
                     merged3_out_5_rest_V => merged_out(5).rest,
                     merged3_out_6_pt_V => merged_out(6).pt,
                     merged3_out_6_eta_V => merged_out(6).eta,
                     merged3_out_6_phi_V => merged_out(6).phi,
                     merged3_out_6_rest_V => merged_out(6).rest,
                     merged3_out_7_pt_V => merged_out(7).pt,
                     merged3_out_7_eta_V => merged_out(7).eta,
                     merged3_out_7_phi_V => merged_out(7).phi,
                     merged3_out_7_rest_V => merged_out(7).rest,
                     merged3_out_8_pt_V => merged_out(8).pt,
                     merged3_out_8_eta_V => merged_out(8).eta,
                     merged3_out_8_phi_V => merged_out(8).phi,
                     merged3_out_8_rest_V => merged_out(8).rest,
                     merged3_out_valid_0 => merged_out_valid(0),
                     merged3_out_valid_1 => merged_out_valid(1),
                     merged3_out_valid_2 => merged_out_valid(2),
                     merged3_out_valid_3 => merged_out_valid(3),
                     merged3_out_valid_4 => merged_out_valid(4),
                     merged3_out_valid_5 => merged_out_valid(5),
                     merged3_out_valid_6 => merged_out_valid(6),
                     merged3_out_valid_7 => merged_out_valid(7),
                     merged3_out_valid_8 => merged_out_valid(8),
                     merged3_out_roll_0 => merged_out_roll(0),
                     merged3_out_roll_1 => merged_out_roll(1),
                     merged3_out_roll_2 => merged_out_roll(2),
                     merged3_out_roll_3 => merged_out_roll(3),
                     merged3_out_roll_4 => merged_out_roll(4),
                     merged3_out_roll_5 => merged_out_roll(5),
                     merged3_out_roll_6 => merged_out_roll(6),
                     merged3_out_roll_7 => merged_out_roll(7),
                     merged3_out_roll_8 => merged_out_roll(8),
                     tracks_out_0_pt_V => tracks_out_0_pt_V,
                     tracks_out_0_eta_V => tracks_out_0_eta_V,
                     tracks_out_0_phi_V => tracks_out_0_phi_V,
                     tracks_out_0_rest_V => tracks_out_0_rest_V,
                     tracks_out_1_eta_V => tracks_out_1_eta_V,
                     tracks_out_1_phi_V => tracks_out_1_phi_V,
                     tracks_out_1_pt_V => tracks_out_1_pt_V,
                     tracks_out_1_rest_V => tracks_out_1_rest_V,
                     tracks_out_2_eta_V => tracks_out_2_eta_V,
                     tracks_out_2_phi_V => tracks_out_2_phi_V,
                     tracks_out_2_pt_V => tracks_out_2_pt_V,
                     tracks_out_2_rest_V => tracks_out_2_rest_V,
                     tracks_out_3_pt_V => tracks_out_3_pt_V,
                     tracks_out_3_eta_V => tracks_out_3_eta_V,
                     tracks_out_3_phi_V => tracks_out_3_phi_V,
                     tracks_out_3_rest_V => tracks_out_3_rest_V,
                     tracks_out_4_eta_V => tracks_out_4_eta_V,
                     tracks_out_4_phi_V => tracks_out_4_phi_V,
                     tracks_out_4_pt_V => tracks_out_4_pt_V,
                     tracks_out_4_rest_V => tracks_out_4_rest_V,
                     tracks_out_5_eta_V => tracks_out_5_eta_V,
                     tracks_out_5_phi_V => tracks_out_5_phi_V,
                     tracks_out_5_pt_V => tracks_out_5_pt_V,
                     tracks_out_5_rest_V => tracks_out_5_rest_V,
                     tracks_out_6_pt_V => tracks_out_6_pt_V,
                     tracks_out_6_eta_V => tracks_out_6_eta_V,
                     tracks_out_6_phi_V => tracks_out_6_phi_V,
                     tracks_out_6_rest_V => tracks_out_6_rest_V,
                     tracks_out_7_eta_V => tracks_out_7_eta_V,
                     tracks_out_7_phi_V => tracks_out_7_phi_V,
                     tracks_out_7_pt_V => tracks_out_7_pt_V,
                     tracks_out_7_rest_V => tracks_out_7_rest_V,
                     tracks_out_8_eta_V => tracks_out_8_eta_V,
                     tracks_out_8_phi_V => tracks_out_8_phi_V,
                     tracks_out_8_pt_V => tracks_out_8_pt_V,
                     tracks_out_8_rest_V => tracks_out_8_rest_V,
                     newevent_out => newevent_out 
                 );


end Behavioral;
